magic
tech sky130A
timestamp 1759050090
<< error_p >>
rect 101 101644 106 101645
rect 124 101644 129 101645
rect 96 101639 134 101640
rect 96 101635 101 101639
rect 128 101635 134 101639
rect 128 101612 129 101635
rect 7921 101508 7926 101509
rect 7944 101508 7949 101509
rect 7916 101503 7954 101504
rect 7916 101499 7921 101503
rect 7948 101499 7954 101503
rect 7948 101476 7949 101499
rect 607 99060 612 99061
rect 630 99060 635 99061
rect 602 99055 640 99056
rect 602 99051 607 99055
rect 634 99051 640 99055
rect 634 99028 635 99051
rect 423 98788 428 98789
rect 446 98788 451 98789
rect 418 98783 456 98784
rect 418 98779 423 98783
rect 450 98779 456 98783
rect 450 98756 451 98779
rect 285 98516 290 98517
rect 308 98516 313 98517
rect 280 98511 318 98512
rect 280 98507 285 98511
rect 312 98507 318 98511
rect 312 98484 313 98507
<< error_s >>
rect 10405 101780 10410 101781
rect 10428 101780 10433 101781
rect 10400 101775 10438 101776
rect 10400 101771 10405 101775
rect 10432 101771 10438 101775
rect 10432 101748 10433 101771
rect 9807 101372 9812 101373
rect 9830 101372 9835 101373
rect 9802 101367 9840 101368
rect 9802 101363 9807 101367
rect 9834 101363 9840 101367
rect 9834 101340 9835 101363
rect 10267 101236 10272 101237
rect 10290 101236 10295 101237
rect 10262 101231 10300 101232
rect 10262 101227 10267 101231
rect 10294 101227 10300 101231
rect 10294 101204 10295 101227
rect 10272 101124 10276 101125
rect 10255 101107 10259 101108
rect 11003 101100 11008 101101
rect 11026 101100 11031 101101
rect 10998 101095 11036 101096
rect 10998 101091 11003 101095
rect 11030 101091 11036 101095
rect 11030 101068 11031 101091
rect 10104 101056 10105 101057
rect 10502 101056 10519 101057
rect 10121 101039 10122 101040
rect 10485 101039 10513 101040
rect 10530 101039 10536 101057
rect 10359 100964 10364 100965
rect 10382 100964 10387 100965
rect 10354 100959 10392 100960
rect 10354 100955 10359 100959
rect 10386 100955 10392 100959
rect 10386 100932 10387 100955
rect 10451 100828 10456 100829
rect 10474 100828 10479 100829
rect 10446 100823 10484 100824
rect 10446 100819 10451 100823
rect 10478 100819 10484 100823
rect 10478 100796 10479 100819
rect 10686 100818 10687 100829
rect 10669 100801 10670 100812
rect 10083 100692 10088 100693
rect 10106 100692 10111 100693
rect 10078 100687 10116 100688
rect 10078 100683 10083 100687
rect 10110 100683 10116 100687
rect 10110 100660 10111 100683
rect 10676 100665 10710 100666
rect 10659 100648 10727 100649
rect 10659 100631 10727 100632
rect 10676 100614 10710 100615
rect 10037 100556 10042 100557
rect 10060 100556 10065 100557
rect 10032 100551 10070 100552
rect 10032 100547 10037 100551
rect 10064 100547 10070 100551
rect 10064 100524 10065 100547
rect 10104 100512 10105 100513
rect 10870 100512 10887 100513
rect 10121 100495 10122 100496
rect 10853 100495 10881 100496
rect 10898 100495 10904 100513
rect 10819 100420 10824 100421
rect 10842 100420 10847 100421
rect 10814 100415 10852 100416
rect 10814 100411 10819 100415
rect 10846 100411 10852 100415
rect 10846 100388 10847 100411
rect 10543 100352 10548 100353
rect 10566 100352 10571 100353
rect 10538 100347 10576 100348
rect 10538 100343 10543 100347
rect 10570 100346 10576 100347
rect 10571 100343 10576 100346
rect 10570 100320 10571 100322
rect 10359 100284 10364 100285
rect 10382 100284 10387 100285
rect 10354 100279 10392 100280
rect 10354 100275 10359 100279
rect 10386 100275 10392 100279
rect 10386 100252 10387 100275
rect 10221 100148 10226 100149
rect 10244 100148 10249 100149
rect 10216 100143 10254 100144
rect 10216 100139 10221 100143
rect 10248 100139 10254 100143
rect 10248 100116 10249 100139
rect 10676 100121 10710 100122
rect 10659 100104 10727 100105
rect 10659 100087 10727 100088
rect 11027 100087 11040 100088
rect 10676 100070 10710 100071
rect 11044 100070 11057 100071
rect 10175 100012 10180 100013
rect 10198 100012 10203 100013
rect 10865 100012 10870 100013
rect 10888 100012 10893 100013
rect 10170 100007 10208 100008
rect 10170 100003 10175 100007
rect 10202 100003 10208 100007
rect 10860 100007 10898 100008
rect 10860 100003 10865 100007
rect 10892 100003 10898 100007
rect 10202 99980 10203 100003
rect 10892 99980 10893 100003
rect 10104 99968 10105 99969
rect 10121 99951 10122 99952
rect 10911 99876 10916 99877
rect 10934 99876 10939 99877
rect 10906 99871 10944 99872
rect 10906 99867 10911 99871
rect 10938 99867 10944 99871
rect 10938 99844 10939 99867
rect 10865 99740 10870 99741
rect 10888 99740 10893 99741
rect 10860 99735 10898 99736
rect 10860 99731 10865 99735
rect 10892 99731 10898 99735
rect 10892 99708 10893 99731
rect 10451 99604 10456 99605
rect 10474 99604 10479 99605
rect 10446 99599 10484 99600
rect 10446 99595 10451 99599
rect 10478 99595 10484 99599
rect 10478 99572 10479 99595
rect 10676 99577 10710 99578
rect 10659 99560 10727 99561
rect 10659 99543 10718 99544
rect 10676 99526 10710 99527
rect 10272 99492 10276 99493
rect 10255 99475 10259 99476
rect 10313 99468 10318 99469
rect 10336 99468 10341 99469
rect 10308 99463 10346 99464
rect 10308 99459 10313 99463
rect 10340 99459 10346 99463
rect 10340 99436 10341 99459
rect 10180 99424 10197 99425
rect 10163 99407 10191 99408
rect 10208 99407 10214 99425
rect 10794 99424 10795 99425
rect 10811 99407 10812 99408
rect 9761 99332 9762 99333
rect 9788 99332 9789 99333
rect 9756 99327 9794 99328
rect 9756 99323 9761 99327
rect 9788 99323 9794 99327
rect 9788 99300 9789 99323
rect 10267 99196 10272 99197
rect 10290 99196 10295 99197
rect 10262 99191 10300 99192
rect 10262 99187 10267 99191
rect 10294 99187 10300 99191
rect 10294 99164 10295 99187
rect 10676 99033 10689 99034
rect 10659 99016 10672 99017
rect 9715 98924 9720 98925
rect 9738 98924 9743 98925
rect 9710 98919 9748 98920
rect 9710 98915 9715 98919
rect 9742 98915 9748 98919
rect 9742 98892 9743 98915
rect 10426 98880 10427 98881
rect 10443 98863 10444 98864
rect 10405 98652 10410 98653
rect 10428 98652 10433 98653
rect 10400 98647 10438 98648
rect 10400 98643 10405 98647
rect 10432 98643 10438 98647
rect 10432 98620 10433 98643
rect 10497 98380 10502 98381
rect 10520 98380 10525 98381
rect 10492 98375 10530 98376
rect 10492 98371 10497 98375
rect 10524 98371 10530 98375
rect 10524 98348 10525 98371
rect 10502 98336 10519 98337
rect 10485 98319 10513 98320
rect 10530 98319 10536 98337
<< locali >>
rect 9720 99305 9737 100580
rect 9766 99339 9783 100478
rect 9812 100155 9829 100750
rect 9858 99509 9875 101056
rect 9950 100767 9967 100954
rect 9783 99322 9784 99331
rect 9766 99306 9784 99322
rect 9766 99169 9783 99306
rect 9904 98591 9921 100410
rect 9950 99951 9967 100274
rect 9950 99679 9967 99866
rect 11100 99407 11117 99730
<< viali >>
rect 10456 101328 10473 101345
rect 10502 101294 10519 101311
rect 10640 101260 10657 101277
rect 10272 101124 10289 101141
rect 9858 101056 9875 101073
rect 10088 101056 10105 101073
rect 10502 101056 10519 101073
rect 9812 100750 9829 100767
rect 9720 100580 9737 100597
rect 9720 99288 9737 99305
rect 9766 100478 9783 100495
rect 9812 100138 9829 100155
rect 10134 101022 10151 101039
rect 10456 101022 10473 101039
rect 9950 100954 9967 100971
rect 10640 100954 10657 100971
rect 10686 100818 10703 100835
rect 10134 100784 10151 100801
rect 10594 100784 10611 100801
rect 10824 100784 10841 100801
rect 9950 100750 9967 100767
rect 10088 100750 10105 100767
rect 10502 100750 10519 100767
rect 10778 100750 10795 100767
rect 11008 100716 11025 100733
rect 10272 100682 10289 100699
rect 10410 100682 10427 100699
rect 10686 100682 10703 100699
rect 10088 100512 10105 100529
rect 10502 100512 10519 100529
rect 10870 100512 10887 100529
rect 10134 100478 10151 100495
rect 10410 100478 10427 100495
rect 10824 100478 10841 100495
rect 10594 100444 10611 100461
rect 9858 99492 9875 99509
rect 9904 100410 9921 100427
rect 10318 100410 10335 100427
rect 10686 100410 10703 100427
rect 11008 100410 11025 100427
rect 9766 99322 9783 99339
rect 9766 99152 9783 99169
rect 9950 100274 9967 100291
rect 10134 100240 10151 100257
rect 10410 100240 10427 100257
rect 10502 100240 10519 100257
rect 10594 100240 10611 100257
rect 10824 100240 10841 100257
rect 10180 100206 10197 100223
rect 10778 100206 10795 100223
rect 11008 100172 11025 100189
rect 10272 100138 10289 100155
rect 10686 100138 10703 100155
rect 10410 100036 10427 100053
rect 10686 100036 10703 100053
rect 10778 100036 10795 100053
rect 10088 99968 10105 99985
rect 10502 99968 10519 99985
rect 9950 99934 9967 99951
rect 10134 99934 10151 99951
rect 10870 99934 10887 99951
rect 10962 99934 10979 99951
rect 10594 99900 10611 99917
rect 9950 99866 9967 99883
rect 10318 99866 10335 99883
rect 11054 99866 11071 99883
rect 10686 99764 10703 99781
rect 10594 99730 10611 99747
rect 11100 99730 11117 99747
rect 10134 99696 10151 99713
rect 9950 99662 9967 99679
rect 10088 99662 10105 99679
rect 10502 99662 10519 99679
rect 10272 99594 10289 99611
rect 10410 99594 10427 99611
rect 10686 99594 10703 99611
rect 10272 99492 10289 99509
rect 10410 99492 10427 99509
rect 10686 99492 10703 99509
rect 11008 99458 11025 99475
rect 10180 99424 10197 99441
rect 10778 99424 10795 99441
rect 10134 99390 10151 99407
rect 10502 99390 10519 99407
rect 10594 99390 10611 99407
rect 10824 99390 10841 99407
rect 11100 99390 11117 99407
rect 10686 99220 10703 99237
rect 10594 99186 10611 99203
rect 10410 99152 10427 99169
rect 10502 99118 10519 99135
rect 10640 98914 10657 98931
rect 10410 98880 10427 98897
rect 10456 98846 10473 98863
rect 10456 98608 10473 98625
rect 9904 98574 9921 98591
rect 10410 98574 10427 98591
rect 10594 98506 10611 98523
rect 10640 98370 10657 98387
rect 10502 98336 10519 98353
rect 10456 98302 10473 98319
<< metal1 >>
rect 10449 101324 10452 101350
rect 10478 101324 10481 101350
rect 10495 101290 10498 101316
rect 10524 101290 10527 101316
rect 10634 101277 10663 101280
rect 10634 101260 10640 101277
rect 10657 101276 10663 101277
rect 10771 101276 10774 101282
rect 10657 101262 10774 101276
rect 10657 101260 10663 101262
rect 10634 101257 10663 101260
rect 10771 101256 10774 101262
rect 10800 101256 10803 101282
rect 10265 101120 10268 101146
rect 10294 101120 10297 101146
rect 9852 101073 9881 101076
rect 9852 101056 9858 101073
rect 9875 101072 9881 101073
rect 10082 101073 10111 101076
rect 10082 101072 10088 101073
rect 9875 101058 10088 101072
rect 9875 101056 9881 101058
rect 9852 101053 9881 101056
rect 10082 101056 10088 101058
rect 10105 101056 10111 101073
rect 10082 101053 10111 101056
rect 10496 101073 10525 101076
rect 10496 101056 10502 101073
rect 10519 101072 10525 101073
rect 10541 101072 10544 101078
rect 10519 101058 10544 101072
rect 10519 101056 10525 101058
rect 10496 101053 10525 101056
rect 10541 101052 10544 101058
rect 10570 101052 10573 101078
rect 10128 101039 10157 101042
rect 10128 101022 10134 101039
rect 10151 101022 10157 101039
rect 10128 101019 10157 101022
rect 10136 101004 10150 101019
rect 10357 101018 10360 101044
rect 10386 101038 10389 101044
rect 10450 101039 10479 101042
rect 10450 101038 10456 101039
rect 10386 101024 10456 101038
rect 10386 101018 10389 101024
rect 10450 101022 10456 101024
rect 10473 101038 10479 101039
rect 10863 101038 10866 101044
rect 10473 101024 10866 101038
rect 10473 101022 10479 101024
rect 10450 101019 10479 101022
rect 10863 101018 10866 101024
rect 10892 101018 10895 101044
rect 10587 101004 10590 101010
rect 10136 100990 10590 101004
rect 10587 100984 10590 100990
rect 10616 100984 10619 101010
rect 9944 100971 9973 100974
rect 9944 100954 9950 100971
rect 9967 100970 9973 100971
rect 10634 100971 10663 100974
rect 10634 100970 10640 100971
rect 9967 100956 10640 100970
rect 9967 100954 9973 100956
rect 9944 100951 9973 100954
rect 10634 100954 10640 100956
rect 10657 100954 10663 100971
rect 10634 100951 10663 100954
rect 10680 100835 10709 100838
rect 10680 100834 10686 100835
rect 10136 100820 10686 100834
rect 10136 100804 10150 100820
rect 10680 100818 10686 100820
rect 10703 100818 10709 100835
rect 10680 100815 10709 100818
rect 10128 100801 10157 100804
rect 10128 100784 10134 100801
rect 10151 100784 10157 100801
rect 10128 100781 10157 100784
rect 10587 100780 10590 100806
rect 10616 100780 10619 100806
rect 10725 100780 10728 100806
rect 10754 100800 10757 100806
rect 10818 100801 10847 100804
rect 10818 100800 10824 100801
rect 10754 100786 10824 100800
rect 10754 100780 10757 100786
rect 10818 100784 10824 100786
rect 10841 100784 10847 100801
rect 10818 100781 10847 100784
rect 9805 100746 9808 100772
rect 9834 100746 9837 100772
rect 9944 100767 9973 100770
rect 9944 100750 9950 100767
rect 9967 100766 9973 100767
rect 10082 100767 10111 100770
rect 10082 100766 10088 100767
rect 9967 100752 10088 100766
rect 9967 100750 9973 100752
rect 9944 100747 9973 100750
rect 10082 100750 10088 100752
rect 10105 100750 10111 100767
rect 10082 100747 10111 100750
rect 10173 100746 10176 100772
rect 10202 100766 10205 100772
rect 10496 100767 10525 100770
rect 10496 100766 10502 100767
rect 10202 100752 10502 100766
rect 10202 100746 10205 100752
rect 10496 100750 10502 100752
rect 10519 100750 10525 100767
rect 10496 100747 10525 100750
rect 10679 100746 10682 100772
rect 10708 100766 10711 100772
rect 10772 100767 10801 100770
rect 10772 100766 10778 100767
rect 10708 100752 10778 100766
rect 10708 100746 10711 100752
rect 10772 100750 10778 100752
rect 10795 100750 10801 100767
rect 10772 100747 10801 100750
rect 10219 100712 10222 100738
rect 10248 100732 10251 100738
rect 11002 100733 11031 100736
rect 11002 100732 11008 100733
rect 10248 100718 11008 100732
rect 10248 100712 10251 100718
rect 11002 100716 11008 100718
rect 11025 100716 11031 100733
rect 11002 100713 11031 100716
rect 99 100678 102 100704
rect 128 100698 131 100704
rect 10266 100699 10295 100702
rect 10266 100698 10272 100699
rect 128 100684 10272 100698
rect 128 100678 131 100684
rect 10266 100682 10272 100684
rect 10289 100682 10295 100699
rect 10266 100679 10295 100682
rect 10403 100678 10406 100704
rect 10432 100678 10435 100704
rect 10680 100699 10709 100702
rect 10680 100682 10686 100699
rect 10703 100698 10709 100699
rect 10955 100698 10958 100704
rect 10703 100684 10958 100698
rect 10703 100682 10709 100684
rect 10680 100679 10709 100682
rect 10955 100678 10958 100684
rect 10984 100678 10987 100704
rect 9714 100597 9743 100600
rect 9714 100580 9720 100597
rect 9737 100596 9743 100597
rect 10403 100596 10406 100602
rect 9737 100582 10406 100596
rect 9737 100580 9743 100582
rect 9714 100577 9743 100580
rect 10403 100576 10406 100582
rect 10432 100576 10435 100602
rect 10909 100562 10912 100568
rect 10504 100548 10912 100562
rect 10035 100508 10038 100534
rect 10064 100528 10067 100534
rect 10504 100532 10518 100548
rect 10909 100542 10912 100548
rect 10938 100542 10941 100568
rect 10082 100529 10111 100532
rect 10082 100528 10088 100529
rect 10064 100514 10088 100528
rect 10064 100508 10067 100514
rect 10082 100512 10088 100514
rect 10105 100512 10111 100529
rect 10082 100509 10111 100512
rect 10496 100529 10525 100532
rect 10496 100512 10502 100529
rect 10519 100512 10525 100529
rect 10496 100509 10525 100512
rect 10864 100529 10893 100532
rect 10864 100512 10870 100529
rect 10887 100528 10893 100529
rect 11047 100528 11050 100534
rect 10887 100514 11050 100528
rect 10887 100512 10893 100514
rect 10864 100509 10893 100512
rect 11047 100508 11050 100514
rect 11076 100508 11079 100534
rect 9760 100495 9789 100498
rect 9760 100478 9766 100495
rect 9783 100494 9789 100495
rect 10128 100495 10157 100498
rect 10128 100494 10134 100495
rect 9783 100480 10134 100494
rect 9783 100478 9789 100480
rect 9760 100475 9789 100478
rect 10128 100478 10134 100480
rect 10151 100478 10157 100495
rect 10128 100475 10157 100478
rect 10403 100474 10406 100500
rect 10432 100474 10435 100500
rect 10818 100495 10847 100498
rect 10818 100494 10824 100495
rect 10550 100480 10824 100494
rect 10357 100440 10360 100466
rect 10386 100460 10389 100466
rect 10550 100460 10564 100480
rect 10818 100478 10824 100480
rect 10841 100478 10847 100495
rect 10818 100475 10847 100478
rect 10386 100446 10564 100460
rect 10588 100461 10617 100464
rect 10386 100440 10389 100446
rect 10588 100444 10594 100461
rect 10611 100460 10617 100461
rect 10725 100460 10728 100466
rect 10611 100446 10728 100460
rect 10611 100444 10617 100446
rect 10588 100441 10617 100444
rect 10725 100440 10728 100446
rect 10754 100440 10757 100466
rect 7919 100406 7922 100432
rect 7948 100426 7951 100432
rect 9898 100427 9927 100430
rect 7948 100412 9667 100426
rect 7948 100406 7951 100412
rect 9653 100290 9667 100412
rect 9898 100410 9904 100427
rect 9921 100426 9927 100427
rect 10312 100427 10341 100430
rect 10312 100426 10318 100427
rect 9921 100412 10318 100426
rect 9921 100410 9927 100412
rect 9898 100407 9927 100410
rect 10312 100410 10318 100412
rect 10335 100410 10341 100427
rect 10312 100407 10341 100410
rect 10633 100406 10636 100432
rect 10662 100426 10665 100432
rect 10680 100427 10709 100430
rect 10680 100426 10686 100427
rect 10662 100412 10686 100426
rect 10662 100406 10665 100412
rect 10680 100410 10686 100412
rect 10703 100410 10709 100427
rect 10680 100407 10709 100410
rect 11002 100427 11031 100430
rect 11002 100410 11008 100427
rect 11025 100426 11031 100427
rect 11025 100412 11070 100426
rect 11025 100410 11031 100412
rect 11002 100407 11031 100410
rect 10081 100304 10084 100330
rect 10110 100324 10113 100330
rect 11056 100324 11070 100412
rect 10110 100310 10518 100324
rect 10110 100304 10113 100310
rect 9944 100291 9973 100294
rect 9944 100290 9950 100291
rect 9653 100276 9950 100290
rect 9944 100274 9950 100276
rect 9967 100290 9973 100291
rect 9967 100276 10426 100290
rect 9967 100274 9973 100276
rect 9944 100271 9973 100274
rect 10127 100236 10130 100262
rect 10156 100236 10159 100262
rect 10412 100260 10426 100276
rect 10504 100260 10518 100310
rect 10642 100310 11070 100324
rect 10404 100257 10433 100260
rect 10404 100240 10410 100257
rect 10427 100240 10433 100257
rect 10404 100237 10433 100240
rect 10496 100257 10525 100260
rect 10496 100240 10502 100257
rect 10519 100240 10525 100257
rect 10496 100237 10525 100240
rect 10541 100236 10544 100262
rect 10570 100256 10573 100262
rect 10588 100257 10617 100260
rect 10588 100256 10594 100257
rect 10570 100242 10594 100256
rect 10570 100236 10573 100242
rect 10588 100240 10594 100242
rect 10611 100240 10617 100257
rect 10588 100237 10617 100240
rect 10174 100223 10203 100226
rect 10174 100206 10180 100223
rect 10197 100222 10203 100223
rect 10642 100222 10656 100310
rect 10817 100236 10820 100262
rect 10846 100236 10849 100262
rect 10197 100208 10656 100222
rect 10197 100206 10203 100208
rect 10174 100203 10203 100206
rect 10771 100202 10774 100228
rect 10800 100202 10803 100228
rect 421 100168 424 100194
rect 450 100188 453 100194
rect 11002 100189 11031 100192
rect 11002 100188 11008 100189
rect 450 100174 11008 100188
rect 450 100168 453 100174
rect 11002 100172 11008 100174
rect 11025 100172 11031 100189
rect 11002 100169 11031 100172
rect 9806 100155 9835 100158
rect 9806 100138 9812 100155
rect 9829 100154 9835 100155
rect 10266 100155 10295 100158
rect 10266 100154 10272 100155
rect 9829 100140 10272 100154
rect 9829 100138 9835 100140
rect 9806 100135 9835 100138
rect 10266 100138 10272 100140
rect 10289 100138 10295 100155
rect 10266 100135 10295 100138
rect 10311 100134 10314 100160
rect 10340 100154 10343 100160
rect 10680 100155 10709 100158
rect 10680 100154 10686 100155
rect 10340 100140 10686 100154
rect 10340 100134 10343 100140
rect 10680 100138 10686 100140
rect 10703 100138 10709 100155
rect 10680 100135 10709 100138
rect 10404 100053 10433 100056
rect 10404 100036 10410 100053
rect 10427 100052 10433 100053
rect 10449 100052 10452 100058
rect 10427 100038 10452 100052
rect 10427 100036 10433 100038
rect 10404 100033 10433 100036
rect 10449 100032 10452 100038
rect 10478 100032 10481 100058
rect 10587 100032 10590 100058
rect 10616 100052 10619 100058
rect 10680 100053 10709 100056
rect 10680 100052 10686 100053
rect 10616 100038 10686 100052
rect 10616 100032 10619 100038
rect 10680 100036 10686 100038
rect 10703 100036 10709 100053
rect 10680 100033 10709 100036
rect 10772 100053 10801 100056
rect 10772 100036 10778 100053
rect 10795 100052 10801 100053
rect 10863 100052 10866 100058
rect 10795 100038 10866 100052
rect 10795 100036 10801 100038
rect 10772 100033 10801 100036
rect 10863 100032 10866 100038
rect 10892 100032 10895 100058
rect 10081 99964 10084 99990
rect 10110 99964 10113 99990
rect 10495 99964 10498 99990
rect 10524 99964 10527 99990
rect 9944 99951 9973 99954
rect 9944 99934 9950 99951
rect 9967 99950 9973 99951
rect 10128 99951 10157 99954
rect 10128 99950 10134 99951
rect 9967 99936 10134 99950
rect 9967 99934 9973 99936
rect 9944 99931 9973 99934
rect 10128 99934 10134 99936
rect 10151 99934 10157 99951
rect 10128 99931 10157 99934
rect 10863 99930 10866 99956
rect 10892 99930 10895 99956
rect 10955 99930 10958 99956
rect 10984 99930 10987 99956
rect 10588 99917 10617 99920
rect 10588 99900 10594 99917
rect 10611 99916 10617 99917
rect 10817 99916 10820 99922
rect 10611 99902 10820 99916
rect 10611 99900 10617 99902
rect 10588 99897 10617 99900
rect 10817 99896 10820 99902
rect 10846 99896 10849 99922
rect 9944 99883 9973 99886
rect 9944 99866 9950 99883
rect 9967 99882 9973 99883
rect 10312 99883 10341 99886
rect 10312 99882 10318 99883
rect 9967 99868 10318 99882
rect 9967 99866 9973 99868
rect 9944 99863 9973 99866
rect 10312 99866 10318 99868
rect 10335 99866 10341 99883
rect 10312 99863 10341 99866
rect 10357 99862 10360 99888
rect 10386 99882 10389 99888
rect 10495 99882 10498 99888
rect 10386 99868 10498 99882
rect 10386 99862 10389 99868
rect 10495 99862 10498 99868
rect 10524 99862 10527 99888
rect 11048 99883 11077 99886
rect 11048 99866 11054 99883
rect 11071 99882 11077 99883
rect 11071 99868 11116 99882
rect 11071 99866 11077 99868
rect 11048 99863 11077 99866
rect 10127 99760 10130 99786
rect 10156 99780 10159 99786
rect 10680 99781 10709 99784
rect 10680 99780 10686 99781
rect 10156 99766 10686 99780
rect 10156 99760 10159 99766
rect 10680 99764 10686 99766
rect 10703 99764 10709 99781
rect 10680 99761 10709 99764
rect 11102 99750 11116 99868
rect 10588 99747 10617 99750
rect 10588 99730 10594 99747
rect 10611 99746 10617 99747
rect 11094 99747 11123 99750
rect 11094 99746 11100 99747
rect 10611 99732 11100 99746
rect 10611 99730 10617 99732
rect 10588 99727 10617 99730
rect 11094 99730 11100 99732
rect 11117 99730 11123 99747
rect 11094 99727 11123 99730
rect 10128 99713 10157 99716
rect 10128 99696 10134 99713
rect 10151 99712 10157 99713
rect 10357 99712 10360 99718
rect 10151 99698 10360 99712
rect 10151 99696 10157 99698
rect 10128 99693 10157 99696
rect 10357 99692 10360 99698
rect 10386 99712 10389 99718
rect 10541 99712 10544 99718
rect 10386 99698 10544 99712
rect 10386 99692 10389 99698
rect 10541 99692 10544 99698
rect 10570 99692 10573 99718
rect 9944 99679 9973 99682
rect 9944 99662 9950 99679
rect 9967 99678 9973 99679
rect 10082 99679 10111 99682
rect 10082 99678 10088 99679
rect 9967 99664 10088 99678
rect 9967 99662 9973 99664
rect 9944 99659 9973 99662
rect 10082 99662 10088 99664
rect 10105 99662 10111 99679
rect 10082 99659 10111 99662
rect 10403 99658 10406 99684
rect 10432 99678 10435 99684
rect 10496 99679 10525 99682
rect 10496 99678 10502 99679
rect 10432 99664 10502 99678
rect 10432 99658 10435 99664
rect 10496 99662 10502 99664
rect 10519 99662 10525 99679
rect 10496 99659 10525 99662
rect 10771 99644 10774 99650
rect 10412 99630 10774 99644
rect 10265 99590 10268 99616
rect 10294 99590 10297 99616
rect 10412 99614 10426 99630
rect 10771 99624 10774 99630
rect 10800 99644 10803 99650
rect 11001 99644 11004 99650
rect 10800 99630 11004 99644
rect 10800 99624 10803 99630
rect 11001 99624 11004 99630
rect 11030 99624 11033 99650
rect 10404 99611 10433 99614
rect 10404 99594 10410 99611
rect 10427 99594 10433 99611
rect 10404 99591 10433 99594
rect 10541 99590 10544 99616
rect 10570 99610 10573 99616
rect 10680 99611 10709 99614
rect 10680 99610 10686 99611
rect 10570 99596 10686 99610
rect 10570 99590 10573 99596
rect 10680 99594 10686 99596
rect 10703 99594 10709 99611
rect 10680 99591 10709 99594
rect 9852 99509 9881 99512
rect 9852 99492 9858 99509
rect 9875 99508 9881 99509
rect 10266 99509 10295 99512
rect 10266 99508 10272 99509
rect 9875 99494 10272 99508
rect 9875 99492 9881 99494
rect 9852 99489 9881 99492
rect 10266 99492 10272 99494
rect 10289 99492 10295 99509
rect 10266 99489 10295 99492
rect 10404 99509 10433 99512
rect 10404 99492 10410 99509
rect 10427 99508 10433 99509
rect 10495 99508 10498 99514
rect 10427 99494 10498 99508
rect 10427 99492 10433 99494
rect 10404 99489 10433 99492
rect 10495 99488 10498 99494
rect 10524 99488 10527 99514
rect 10680 99509 10709 99512
rect 10680 99492 10686 99509
rect 10703 99508 10709 99509
rect 10725 99508 10728 99514
rect 10703 99494 10728 99508
rect 10703 99492 10709 99494
rect 10680 99489 10709 99492
rect 10725 99488 10728 99494
rect 10754 99488 10757 99514
rect 283 99454 286 99480
rect 312 99474 315 99480
rect 11002 99475 11031 99478
rect 11002 99474 11008 99475
rect 312 99460 11008 99474
rect 312 99454 315 99460
rect 11002 99458 11008 99460
rect 11025 99458 11031 99475
rect 11002 99455 11031 99458
rect 10173 99420 10176 99446
rect 10202 99420 10205 99446
rect 10633 99420 10636 99446
rect 10662 99440 10665 99446
rect 10772 99441 10801 99444
rect 10772 99440 10778 99441
rect 10662 99426 10778 99440
rect 10662 99420 10665 99426
rect 10772 99424 10778 99426
rect 10795 99424 10801 99441
rect 10772 99421 10801 99424
rect 10128 99407 10157 99410
rect 10128 99390 10134 99407
rect 10151 99390 10157 99407
rect 10128 99387 10157 99390
rect 9759 99318 9762 99344
rect 9788 99318 9791 99344
rect 10136 99338 10150 99387
rect 10495 99386 10498 99412
rect 10524 99386 10527 99412
rect 10541 99386 10544 99412
rect 10570 99406 10573 99412
rect 10588 99407 10617 99410
rect 10588 99406 10594 99407
rect 10570 99392 10594 99406
rect 10570 99386 10573 99392
rect 10588 99390 10594 99392
rect 10611 99390 10617 99407
rect 10588 99387 10617 99390
rect 10818 99407 10847 99410
rect 10818 99390 10824 99407
rect 10841 99406 10847 99407
rect 11094 99407 11123 99410
rect 11094 99406 11100 99407
rect 10841 99392 11100 99406
rect 10841 99390 10847 99392
rect 10818 99387 10847 99390
rect 11094 99390 11100 99392
rect 11117 99390 11123 99407
rect 11094 99387 11123 99390
rect 10504 99372 10518 99386
rect 11001 99372 11004 99378
rect 10504 99358 11004 99372
rect 11001 99352 11004 99358
rect 11030 99352 11033 99378
rect 9998 99324 10150 99338
rect 9713 99284 9716 99310
rect 9742 99304 9745 99310
rect 9998 99304 10012 99324
rect 9742 99290 10012 99304
rect 9742 99284 9745 99290
rect 10357 99216 10360 99242
rect 10386 99236 10389 99242
rect 10680 99237 10709 99240
rect 10680 99236 10686 99237
rect 10386 99222 10686 99236
rect 10386 99216 10389 99222
rect 10680 99220 10686 99222
rect 10703 99220 10709 99237
rect 10680 99217 10709 99220
rect 10587 99182 10590 99208
rect 10616 99182 10619 99208
rect 9760 99169 9789 99172
rect 9760 99152 9766 99169
rect 9783 99168 9789 99169
rect 10404 99169 10433 99172
rect 10404 99168 10410 99169
rect 9783 99154 10410 99168
rect 9783 99152 9789 99154
rect 9760 99149 9789 99152
rect 10404 99152 10410 99154
rect 10427 99152 10433 99169
rect 10404 99149 10433 99152
rect 10035 99114 10038 99140
rect 10064 99134 10067 99140
rect 10496 99135 10525 99138
rect 10496 99134 10502 99135
rect 10064 99120 10502 99134
rect 10064 99114 10067 99120
rect 10496 99118 10502 99120
rect 10519 99118 10525 99135
rect 10496 99115 10525 99118
rect 10633 98910 10636 98936
rect 10662 98910 10665 98936
rect 10403 98876 10406 98902
rect 10432 98876 10435 98902
rect 10450 98863 10479 98866
rect 10450 98846 10456 98863
rect 10473 98862 10479 98863
rect 10771 98862 10774 98868
rect 10473 98848 10774 98862
rect 10473 98846 10479 98848
rect 10450 98843 10479 98846
rect 10771 98842 10774 98848
rect 10800 98842 10803 98868
rect 10587 98692 10590 98698
rect 10458 98678 10590 98692
rect 10458 98628 10472 98678
rect 10587 98672 10590 98678
rect 10616 98672 10619 98698
rect 10450 98625 10479 98628
rect 10450 98608 10456 98625
rect 10473 98608 10479 98625
rect 10450 98605 10479 98608
rect 9898 98591 9927 98594
rect 9898 98574 9904 98591
rect 9921 98590 9927 98591
rect 10404 98591 10433 98594
rect 10404 98590 10410 98591
rect 9921 98576 10410 98590
rect 9921 98574 9927 98576
rect 9898 98571 9927 98574
rect 10404 98574 10410 98576
rect 10427 98574 10433 98591
rect 10404 98571 10433 98574
rect 605 98502 608 98528
rect 634 98522 637 98528
rect 10588 98523 10617 98526
rect 10588 98522 10594 98523
rect 634 98508 10594 98522
rect 634 98502 637 98508
rect 10588 98506 10594 98508
rect 10611 98506 10617 98523
rect 10588 98503 10617 98506
rect 10634 98387 10663 98390
rect 10634 98370 10640 98387
rect 10657 98386 10663 98387
rect 10679 98386 10682 98392
rect 10657 98372 10682 98386
rect 10657 98370 10663 98372
rect 10634 98367 10663 98370
rect 10679 98366 10682 98372
rect 10708 98366 10711 98392
rect 10496 98353 10525 98356
rect 10496 98336 10502 98353
rect 10519 98352 10525 98353
rect 10909 98352 10912 98358
rect 10519 98338 10912 98352
rect 10519 98336 10525 98338
rect 10496 98333 10525 98336
rect 10909 98332 10912 98338
rect 10938 98332 10941 98358
rect 10449 98298 10452 98324
rect 10478 98298 10481 98324
<< via1 >>
rect 10452 101345 10478 101350
rect 10452 101328 10456 101345
rect 10456 101328 10473 101345
rect 10473 101328 10478 101345
rect 10452 101324 10478 101328
rect 10498 101311 10524 101316
rect 10498 101294 10502 101311
rect 10502 101294 10519 101311
rect 10519 101294 10524 101311
rect 10498 101290 10524 101294
rect 10774 101256 10800 101282
rect 10268 101141 10294 101146
rect 10268 101124 10272 101141
rect 10272 101124 10289 101141
rect 10289 101124 10294 101141
rect 10268 101120 10294 101124
rect 10544 101052 10570 101078
rect 10360 101018 10386 101044
rect 10866 101018 10892 101044
rect 10590 100984 10616 101010
rect 10590 100801 10616 100806
rect 10590 100784 10594 100801
rect 10594 100784 10611 100801
rect 10611 100784 10616 100801
rect 10590 100780 10616 100784
rect 10728 100780 10754 100806
rect 9808 100767 9834 100772
rect 9808 100750 9812 100767
rect 9812 100750 9829 100767
rect 9829 100750 9834 100767
rect 9808 100746 9834 100750
rect 10176 100746 10202 100772
rect 10682 100746 10708 100772
rect 10222 100712 10248 100738
rect 102 100678 128 100704
rect 10406 100699 10432 100704
rect 10406 100682 10410 100699
rect 10410 100682 10427 100699
rect 10427 100682 10432 100699
rect 10406 100678 10432 100682
rect 10958 100678 10984 100704
rect 10406 100576 10432 100602
rect 10038 100508 10064 100534
rect 10912 100542 10938 100568
rect 11050 100508 11076 100534
rect 10406 100495 10432 100500
rect 10406 100478 10410 100495
rect 10410 100478 10427 100495
rect 10427 100478 10432 100495
rect 10406 100474 10432 100478
rect 10360 100440 10386 100466
rect 10728 100440 10754 100466
rect 7922 100406 7948 100432
rect 10636 100406 10662 100432
rect 10084 100304 10110 100330
rect 10130 100257 10156 100262
rect 10130 100240 10134 100257
rect 10134 100240 10151 100257
rect 10151 100240 10156 100257
rect 10130 100236 10156 100240
rect 10544 100236 10570 100262
rect 10820 100257 10846 100262
rect 10820 100240 10824 100257
rect 10824 100240 10841 100257
rect 10841 100240 10846 100257
rect 10820 100236 10846 100240
rect 10774 100223 10800 100228
rect 10774 100206 10778 100223
rect 10778 100206 10795 100223
rect 10795 100206 10800 100223
rect 10774 100202 10800 100206
rect 424 100168 450 100194
rect 10314 100134 10340 100160
rect 10452 100032 10478 100058
rect 10590 100032 10616 100058
rect 10866 100032 10892 100058
rect 10084 99985 10110 99990
rect 10084 99968 10088 99985
rect 10088 99968 10105 99985
rect 10105 99968 10110 99985
rect 10084 99964 10110 99968
rect 10498 99985 10524 99990
rect 10498 99968 10502 99985
rect 10502 99968 10519 99985
rect 10519 99968 10524 99985
rect 10498 99964 10524 99968
rect 10866 99951 10892 99956
rect 10866 99934 10870 99951
rect 10870 99934 10887 99951
rect 10887 99934 10892 99951
rect 10866 99930 10892 99934
rect 10958 99951 10984 99956
rect 10958 99934 10962 99951
rect 10962 99934 10979 99951
rect 10979 99934 10984 99951
rect 10958 99930 10984 99934
rect 10820 99896 10846 99922
rect 10360 99862 10386 99888
rect 10498 99862 10524 99888
rect 10130 99760 10156 99786
rect 10360 99692 10386 99718
rect 10544 99692 10570 99718
rect 10406 99658 10432 99684
rect 10268 99611 10294 99616
rect 10268 99594 10272 99611
rect 10272 99594 10289 99611
rect 10289 99594 10294 99611
rect 10268 99590 10294 99594
rect 10774 99624 10800 99650
rect 11004 99624 11030 99650
rect 10544 99590 10570 99616
rect 10498 99488 10524 99514
rect 10728 99488 10754 99514
rect 286 99454 312 99480
rect 10176 99441 10202 99446
rect 10176 99424 10180 99441
rect 10180 99424 10197 99441
rect 10197 99424 10202 99441
rect 10176 99420 10202 99424
rect 10636 99420 10662 99446
rect 9762 99339 9788 99344
rect 9762 99322 9766 99339
rect 9766 99322 9783 99339
rect 9783 99322 9788 99339
rect 9762 99318 9788 99322
rect 10498 99407 10524 99412
rect 10498 99390 10502 99407
rect 10502 99390 10519 99407
rect 10519 99390 10524 99407
rect 10498 99386 10524 99390
rect 10544 99386 10570 99412
rect 11004 99352 11030 99378
rect 9716 99305 9742 99310
rect 9716 99288 9720 99305
rect 9720 99288 9737 99305
rect 9737 99288 9742 99305
rect 9716 99284 9742 99288
rect 10360 99216 10386 99242
rect 10590 99203 10616 99208
rect 10590 99186 10594 99203
rect 10594 99186 10611 99203
rect 10611 99186 10616 99203
rect 10590 99182 10616 99186
rect 10038 99114 10064 99140
rect 10636 98931 10662 98936
rect 10636 98914 10640 98931
rect 10640 98914 10657 98931
rect 10657 98914 10662 98931
rect 10636 98910 10662 98914
rect 10406 98897 10432 98902
rect 10406 98880 10410 98897
rect 10410 98880 10427 98897
rect 10427 98880 10432 98897
rect 10406 98876 10432 98880
rect 10774 98842 10800 98868
rect 10590 98672 10616 98698
rect 608 98502 634 98528
rect 10682 98366 10708 98392
rect 10912 98332 10938 98358
rect 10452 98319 10478 98324
rect 10452 98302 10456 98319
rect 10456 98302 10473 98319
rect 10473 98302 10478 98319
rect 10452 98298 10478 98302
<< metal2 >>
rect 10405 101776 10433 101780
rect 10405 101743 10433 101748
rect 101 101640 129 101644
rect 101 101607 129 101612
rect 108 100707 122 101607
rect 7921 101504 7949 101508
rect 7921 101471 7949 101476
rect 102 100704 128 100707
rect 102 100675 128 100678
rect 7928 100435 7942 101471
rect 10412 101437 10426 101743
rect 10412 101423 10518 101437
rect 9807 101368 9835 101372
rect 9807 101335 9835 101340
rect 10452 101350 10478 101353
rect 9814 100775 9828 101335
rect 10452 101321 10478 101324
rect 10267 101232 10295 101236
rect 10267 101199 10295 101204
rect 10274 101149 10288 101199
rect 10268 101146 10294 101149
rect 10268 101117 10294 101120
rect 10360 101044 10386 101047
rect 10360 101015 10386 101018
rect 10366 100964 10380 101015
rect 10359 100960 10387 100964
rect 10359 100927 10387 100932
rect 10458 100828 10472 101321
rect 10504 101319 10518 101423
rect 10498 101316 10524 101319
rect 10498 101287 10524 101290
rect 10451 100824 10479 100828
rect 10451 100791 10479 100796
rect 9808 100772 9834 100775
rect 9808 100743 9834 100746
rect 10176 100772 10202 100775
rect 10176 100743 10202 100746
rect 10083 100688 10111 100692
rect 10083 100655 10111 100660
rect 10037 100552 10065 100556
rect 10037 100519 10038 100524
rect 10064 100519 10065 100524
rect 10038 100505 10064 100508
rect 7922 100432 7948 100435
rect 7922 100403 7948 100406
rect 424 100194 450 100197
rect 424 100165 450 100168
rect 286 99480 312 99483
rect 286 99451 312 99454
rect 292 98516 306 99451
rect 430 98788 444 100165
rect 9762 99344 9788 99347
rect 9761 99328 9762 99332
rect 9788 99328 9789 99332
rect 9716 99310 9742 99313
rect 9761 99295 9789 99300
rect 9716 99281 9742 99284
rect 607 99056 635 99060
rect 607 99023 635 99028
rect 423 98784 451 98788
rect 423 98751 451 98756
rect 614 98531 628 99023
rect 9722 98924 9736 99281
rect 10044 99143 10058 100505
rect 10090 100333 10104 100655
rect 10084 100330 10110 100333
rect 10084 100301 10110 100304
rect 10090 99993 10104 100301
rect 10130 100262 10156 100265
rect 10130 100233 10156 100236
rect 10084 99990 10110 99993
rect 10084 99961 10110 99964
rect 10136 99789 10150 100233
rect 10182 100012 10196 100743
rect 10222 100738 10248 100741
rect 10222 100709 10248 100712
rect 10228 100148 10242 100709
rect 10406 100704 10432 100707
rect 10406 100675 10432 100678
rect 10412 100605 10426 100675
rect 10406 100602 10432 100605
rect 10406 100573 10432 100576
rect 10406 100500 10432 100503
rect 10406 100471 10432 100474
rect 10360 100466 10386 100469
rect 10360 100437 10386 100440
rect 10366 100284 10380 100437
rect 10359 100280 10387 100284
rect 10359 100247 10387 100252
rect 10314 100160 10340 100163
rect 10221 100144 10249 100148
rect 10314 100131 10340 100134
rect 10221 100111 10249 100116
rect 10175 100008 10203 100012
rect 10175 99975 10203 99980
rect 10130 99786 10156 99789
rect 10130 99757 10156 99760
rect 10182 99449 10196 99975
rect 10268 99616 10294 99619
rect 10268 99587 10294 99590
rect 10176 99446 10202 99449
rect 10176 99417 10202 99420
rect 10274 99196 10288 99587
rect 10320 99468 10334 100131
rect 10366 99891 10380 100247
rect 10360 99888 10386 99891
rect 10360 99859 10386 99862
rect 10412 99729 10426 100471
rect 10458 100061 10472 100791
rect 10452 100058 10478 100061
rect 10452 100029 10478 100032
rect 10504 99993 10518 101287
rect 10774 101282 10800 101285
rect 10774 101253 10800 101256
rect 10544 101078 10570 101081
rect 10544 101049 10570 101052
rect 10550 100352 10564 101049
rect 10590 101010 10616 101013
rect 10590 100981 10616 100984
rect 10596 100809 10610 100981
rect 10590 100806 10616 100809
rect 10590 100777 10616 100780
rect 10728 100806 10754 100809
rect 10728 100777 10754 100780
rect 10543 100348 10571 100352
rect 10543 100315 10571 100320
rect 10544 100262 10570 100265
rect 10544 100233 10570 100236
rect 10498 99990 10524 99993
rect 10498 99961 10524 99964
rect 10498 99888 10524 99891
rect 10498 99859 10524 99862
rect 10360 99718 10386 99721
rect 10412 99715 10472 99729
rect 10360 99689 10386 99692
rect 10313 99464 10341 99468
rect 10313 99431 10341 99436
rect 10366 99245 10380 99689
rect 10406 99684 10432 99687
rect 10406 99655 10432 99658
rect 10360 99242 10386 99245
rect 10360 99213 10386 99216
rect 10267 99192 10295 99196
rect 10267 99159 10295 99164
rect 10038 99140 10064 99143
rect 10038 99111 10064 99114
rect 9715 98920 9743 98924
rect 10412 98905 10426 99655
rect 10458 99604 10472 99715
rect 10451 99600 10479 99604
rect 10451 99567 10479 99572
rect 9715 98887 9743 98892
rect 10406 98902 10432 98905
rect 10406 98873 10432 98876
rect 10412 98652 10426 98873
rect 10405 98648 10433 98652
rect 10405 98615 10433 98620
rect 608 98528 634 98531
rect 285 98512 313 98516
rect 608 98499 634 98502
rect 285 98479 313 98484
rect 10458 98327 10472 99567
rect 10504 99517 10518 99859
rect 10550 99721 10564 100233
rect 10596 100061 10610 100777
rect 10682 100772 10708 100775
rect 10682 100743 10708 100746
rect 10636 100432 10662 100435
rect 10636 100403 10662 100406
rect 10590 100058 10616 100061
rect 10590 100029 10616 100032
rect 10544 99718 10570 99721
rect 10544 99689 10570 99692
rect 10544 99616 10570 99619
rect 10544 99587 10570 99590
rect 10498 99514 10524 99517
rect 10498 99485 10524 99488
rect 10550 99415 10564 99587
rect 10642 99525 10656 100403
rect 10596 99511 10656 99525
rect 10498 99412 10524 99415
rect 10498 99383 10524 99386
rect 10544 99412 10570 99415
rect 10544 99383 10570 99386
rect 10504 98380 10518 99383
rect 10596 99211 10610 99511
rect 10636 99446 10662 99449
rect 10636 99417 10662 99420
rect 10590 99208 10616 99211
rect 10590 99179 10616 99182
rect 10596 98701 10610 99179
rect 10642 98939 10656 99417
rect 10636 98936 10662 98939
rect 10636 98907 10662 98910
rect 10590 98698 10616 98701
rect 10590 98669 10616 98672
rect 10688 98395 10702 100743
rect 10734 100469 10748 100777
rect 10728 100466 10754 100469
rect 10728 100437 10754 100440
rect 10734 99517 10748 100437
rect 10780 100231 10794 101253
rect 11003 101096 11031 101100
rect 11003 101063 11031 101068
rect 10866 101044 10892 101047
rect 10866 101015 10892 101018
rect 10819 100416 10847 100420
rect 10819 100383 10847 100388
rect 10826 100265 10840 100383
rect 10820 100262 10846 100265
rect 10820 100233 10846 100236
rect 10774 100228 10800 100231
rect 10774 100199 10800 100202
rect 10826 99925 10840 100233
rect 10872 100061 10886 101015
rect 10958 100704 10984 100707
rect 10958 100675 10984 100678
rect 10912 100568 10938 100571
rect 10912 100539 10938 100542
rect 10866 100058 10892 100061
rect 10866 100029 10892 100032
rect 10865 100008 10893 100012
rect 10865 99975 10893 99980
rect 10872 99959 10886 99975
rect 10866 99956 10892 99959
rect 10866 99927 10892 99930
rect 10820 99922 10846 99925
rect 10820 99893 10846 99896
rect 10872 99740 10886 99927
rect 10918 99876 10932 100539
rect 10964 99959 10978 100675
rect 10958 99956 10984 99959
rect 10958 99927 10984 99930
rect 10911 99872 10939 99876
rect 10911 99839 10939 99844
rect 10865 99736 10893 99740
rect 10865 99703 10893 99708
rect 10774 99650 10800 99653
rect 10774 99621 10800 99624
rect 10728 99514 10754 99517
rect 10728 99485 10754 99488
rect 10780 98871 10794 99621
rect 10774 98868 10800 98871
rect 10774 98839 10800 98842
rect 10682 98392 10708 98395
rect 10497 98376 10525 98380
rect 10682 98363 10708 98366
rect 10918 98361 10932 99839
rect 11010 99653 11024 101063
rect 11050 100534 11076 100537
rect 11050 100505 11076 100508
rect 11004 99650 11030 99653
rect 11004 99621 11030 99624
rect 11056 99593 11070 100505
rect 11010 99579 11070 99593
rect 11010 99381 11024 99579
rect 11004 99378 11030 99381
rect 11004 99349 11030 99352
rect 10497 98343 10525 98348
rect 10912 98358 10938 98361
rect 10912 98329 10938 98332
rect 10452 98324 10478 98327
rect 10452 98295 10478 98298
<< via2 >>
rect 10405 101748 10433 101776
rect 101 101612 129 101640
rect 7921 101476 7949 101504
rect 9807 101340 9835 101368
rect 10267 101204 10295 101232
rect 10359 100932 10387 100960
rect 10451 100796 10479 100824
rect 10083 100660 10111 100688
rect 10037 100534 10065 100552
rect 10037 100524 10038 100534
rect 10038 100524 10064 100534
rect 10064 100524 10065 100534
rect 9761 99318 9762 99328
rect 9762 99318 9788 99328
rect 9788 99318 9789 99328
rect 9761 99300 9789 99318
rect 607 99028 635 99056
rect 423 98756 451 98784
rect 10359 100252 10387 100280
rect 10221 100116 10249 100144
rect 10175 99980 10203 100008
rect 10543 100320 10571 100348
rect 10313 99436 10341 99464
rect 10267 99164 10295 99192
rect 9715 98892 9743 98920
rect 10451 99572 10479 99600
rect 10405 98620 10433 98648
rect 285 98484 313 98512
rect 11003 101068 11031 101096
rect 10819 100388 10847 100416
rect 10865 99980 10893 100008
rect 10911 99844 10939 99872
rect 10865 99708 10893 99736
rect 10497 98348 10525 98376
<< metal3 >>
rect 10402 101777 10435 101778
rect 0 101776 10435 101777
rect 0 101748 10405 101776
rect 10433 101748 10435 101776
rect 0 101747 10435 101748
rect 10402 101745 10435 101747
rect 98 101641 131 101642
rect 0 101640 131 101641
rect 0 101612 101 101640
rect 129 101612 131 101640
rect 0 101611 131 101612
rect 98 101609 131 101611
rect 7918 101505 7951 101506
rect 0 101504 7951 101505
rect 0 101476 7921 101504
rect 7949 101476 7951 101504
rect 0 101475 7951 101476
rect 7918 101473 7951 101475
rect 9804 101369 9837 101370
rect 0 101368 9837 101369
rect 0 101340 9807 101368
rect 9835 101340 9837 101368
rect 0 101339 9837 101340
rect 9804 101337 9837 101339
rect 10264 101233 10297 101234
rect 0 101232 10297 101233
rect 0 101204 10267 101232
rect 10295 101204 10297 101232
rect 0 101203 10297 101204
rect 10264 101201 10297 101203
rect 11000 101097 11033 101098
rect 0 101096 11033 101097
rect 0 101068 11003 101096
rect 11031 101068 11033 101096
rect 0 101067 11033 101068
rect 11000 101065 11033 101067
rect 10356 100961 10389 100962
rect 0 100960 10389 100961
rect 0 100932 10359 100960
rect 10387 100932 10389 100960
rect 0 100931 10389 100932
rect 10356 100929 10389 100931
rect 10448 100825 10481 100826
rect 0 100824 10481 100825
rect 0 100796 10451 100824
rect 10479 100796 10481 100824
rect 0 100795 10481 100796
rect 10448 100793 10481 100795
rect 10080 100689 10113 100690
rect 0 100688 10113 100689
rect 0 100660 10083 100688
rect 10111 100660 10113 100688
rect 0 100659 10113 100660
rect 10080 100657 10113 100659
rect 10034 100553 10067 100554
rect 0 100552 10067 100553
rect 0 100524 10037 100552
rect 10065 100524 10067 100552
rect 0 100523 10067 100524
rect 10034 100521 10067 100523
rect 10816 100417 10849 100418
rect 0 100416 10849 100417
rect 0 100388 10819 100416
rect 10847 100388 10849 100416
rect 0 100387 10849 100388
rect 10816 100385 10849 100387
rect 10540 100349 10573 100350
rect 10540 100348 10641 100349
rect 10540 100320 10543 100348
rect 10571 100320 10641 100348
rect 10540 100319 10641 100320
rect 10540 100317 10573 100319
rect 10356 100281 10389 100282
rect 0 100280 10389 100281
rect 0 100252 10359 100280
rect 10387 100252 10389 100280
rect 0 100251 10389 100252
rect 10356 100249 10389 100251
rect 10218 100145 10251 100146
rect 0 100144 10251 100145
rect 0 100116 10221 100144
rect 10249 100116 10251 100144
rect 0 100115 10251 100116
rect 10218 100113 10251 100115
rect 10172 100009 10205 100010
rect 0 100008 10205 100009
rect 0 99980 10175 100008
rect 10203 99980 10205 100008
rect 0 99979 10205 99980
rect 10611 100009 10641 100319
rect 10862 100009 10895 100010
rect 10611 100008 10895 100009
rect 10611 99980 10865 100008
rect 10893 99980 10895 100008
rect 10611 99979 10895 99980
rect 10172 99977 10205 99979
rect 10862 99977 10895 99979
rect 10908 99873 10941 99874
rect 0 99872 10941 99873
rect 0 99844 10911 99872
rect 10939 99844 10941 99872
rect 0 99843 10941 99844
rect 10908 99841 10941 99843
rect 10862 99737 10895 99738
rect 0 99736 10895 99737
rect 0 99708 10865 99736
rect 10893 99708 10895 99736
rect 0 99707 10895 99708
rect 10862 99705 10895 99707
rect 10448 99601 10481 99602
rect 0 99600 10481 99601
rect 0 99572 10451 99600
rect 10479 99572 10481 99600
rect 0 99571 10481 99572
rect 10448 99569 10481 99571
rect 10310 99465 10343 99466
rect 0 99464 10343 99465
rect 0 99436 10313 99464
rect 10341 99436 10343 99464
rect 0 99435 10343 99436
rect 10310 99433 10343 99435
rect 9758 99329 9791 99330
rect 0 99328 9791 99329
rect 0 99300 9761 99328
rect 9789 99300 9791 99328
rect 0 99299 9791 99300
rect 9758 99297 9791 99299
rect 10264 99193 10297 99194
rect 0 99192 10297 99193
rect 0 99164 10267 99192
rect 10295 99164 10297 99192
rect 0 99163 10297 99164
rect 10264 99161 10297 99163
rect 604 99057 637 99058
rect 0 99056 637 99057
rect 0 99028 607 99056
rect 635 99028 637 99056
rect 0 99027 637 99028
rect 604 99025 637 99027
rect 9712 98921 9745 98922
rect 0 98920 9745 98921
rect 0 98892 9715 98920
rect 9743 98892 9745 98920
rect 0 98891 9745 98892
rect 9712 98889 9745 98891
rect 420 98785 453 98786
rect 0 98784 453 98785
rect 0 98756 423 98784
rect 451 98756 453 98784
rect 0 98755 453 98756
rect 420 98753 453 98755
rect 10402 98649 10435 98650
rect 0 98648 10435 98649
rect 0 98620 10405 98648
rect 10433 98620 10435 98648
rect 0 98619 10435 98620
rect 10402 98617 10435 98619
rect 282 98513 315 98514
rect 0 98512 315 98513
rect 0 98484 285 98512
rect 313 98484 315 98512
rect 0 98483 315 98484
rect 282 98481 315 98483
rect 10494 98377 10527 98378
rect 0 98376 10527 98377
rect 0 98348 10497 98376
rect 10525 98348 10527 98376
rect 0 98347 10527 98348
rect 10494 98345 10527 98347
<< metal4 >>
rect 215 0 245 80
rect 399 0 429 80
use sky130_fd_sc_hd__xnor2_1  UUT_C1__07_
timestamp 1759050090
transform 1 0 10350 0 -1 101456
box -19 -24 341 296
use sky130_fd_sc_hd__maj3_1  UUT_C1__08_
timestamp 1759050090
transform 1 0 10350 0 1 99824
box -19 -24 387 296
use sky130_fd_sc_hd__xnor2_1  UUT_C1__09_
timestamp 1759050090
transform 1 0 10028 0 1 99280
box -19 -24 341 296
use sky130_fd_sc_hd__maj3_1  UUT_C1__10_
timestamp 1759050090
transform 1 0 10350 0 -1 100912
box -19 -24 387 296
use sky130_fd_sc_hd__xnor2_1  UUT_C1__11_
timestamp 1759050090
transform 1 0 10350 0 1 100912
box -19 -24 341 296
use sky130_fd_sc_hd__maj3_1  UUT_C1__12_
timestamp 1759050090
transform 1 0 10718 0 1 99824
box -19 -24 387 296
use sky130_fd_sc_hd__xnor2_1  UUT_C1__13_
timestamp 1759050090
transform 1 0 10350 0 1 98736
box -19 -24 341 296
use sky130_fd_sc_hd__maj3_1  UUT_C1__14_
timestamp 1759050090
transform 1 0 10350 0 -1 99824
box -19 -24 387 296
use sky130_fd_sc_hd__xnor2_1  UUT_C1__15_
timestamp 1759050090
transform 1 0 10718 0 -1 100368
box -19 -24 341 296
use sky130_fd_sc_hd__xnor2_1  UUT_C1__16_
timestamp 1759050090
transform 1 0 10028 0 1 100912
box -19 -24 341 296
use sky130_fd_sc_hd__xnor2_1  UUT_C1__17_
timestamp 1759050090
transform 1 0 10028 0 -1 100912
box -19 -24 341 296
use sky130_fd_sc_hd__xnor2_1  UUT_C1__18_
timestamp 1759050090
transform 1 0 10718 0 1 99280
box -19 -24 341 296
use sky130_fd_sc_hd__xnor2_1  UUT_C2__07_
timestamp 1759050090
transform 1 0 10718 0 1 100368
box -19 -24 341 296
use sky130_fd_sc_hd__maj3_1  UUT_C2__08_
timestamp 1759050090
transform 1 0 10350 0 1 99280
box -19 -24 387 296
use sky130_fd_sc_hd__xnor2_1  UUT_C2__09_
timestamp 1759050090
transform 1 0 10350 0 1 98192
box -19 -24 341 296
use sky130_fd_sc_hd__maj3_1  UUT_C2__10_
timestamp 1759050090
transform 1 0 10350 0 1 100368
box -19 -24 387 296
use sky130_fd_sc_hd__xnor2_1  UUT_C2__11_
timestamp 1759050090
transform 1 0 10028 0 1 100368
box -19 -24 341 296
use sky130_fd_sc_hd__maj3_1  UUT_C2__12_
timestamp 1759050090
transform 1 0 10350 0 -1 99280
box -19 -24 387 296
use sky130_fd_sc_hd__xnor2_1  UUT_C2__13_
timestamp 1759050090
transform 1 0 10028 0 1 99824
box -19 -24 341 296
use sky130_fd_sc_hd__maj3_1  UUT_C2__14_
timestamp 1759050090
transform 1 0 10350 0 -1 100368
box -19 -24 387 296
use sky130_fd_sc_hd__xnor2_1  UUT_C2__15_
timestamp 1759050090
transform 1 0 10028 0 -1 100368
box -19 -24 341 296
use sky130_fd_sc_hd__xnor2_1  UUT_C2__16_
timestamp 1759050090
transform 1 0 10718 0 -1 100912
box -19 -24 341 296
use sky130_fd_sc_hd__xnor2_1  UUT_C2__17_
timestamp 1759050090
transform 1 0 10350 0 -1 98736
box -19 -24 341 296
use sky130_fd_sc_hd__xnor2_1  UUT_C2__18_
timestamp 1759050090
transform 1 0 10028 0 -1 99824
box -19 -24 341 296
<< labels >>
flabel metal3 s 0 101747 80 101777 0 FreeSans 240 0 0 0 A[0]
port 0 nsew signal input
flabel metal3 s 0 99979 80 100009 0 FreeSans 240 0 0 0 A[1]
port 1 nsew signal input
flabel metal3 s 0 99707 80 99737 0 FreeSans 240 0 0 0 A[2]
port 2 nsew signal input
flabel metal3 s 0 98619 80 98649 0 FreeSans 240 0 0 0 A[3]
port 3 nsew signal input
flabel metal3 s 0 98347 80 98377 0 FreeSans 240 0 0 0 A[4]
port 4 nsew signal input
flabel metal3 s 0 99843 80 99873 0 FreeSans 240 0 0 0 A[5]
port 5 nsew signal input
flabel metal3 s 0 100523 80 100553 0 FreeSans 240 0 0 0 A[6]
port 6 nsew signal input
flabel metal3 s 0 100659 80 100689 0 FreeSans 240 0 0 0 A[7]
port 7 nsew signal input
flabel metal3 s 0 100795 80 100825 0 FreeSans 240 0 0 0 B[0]
port 8 nsew signal input
flabel metal3 s 0 98891 80 98921 0 FreeSans 240 0 0 0 B[1]
port 9 nsew signal input
flabel metal3 s 0 100931 80 100961 0 FreeSans 240 0 0 0 B[2]
port 10 nsew signal input
flabel metal3 s 0 101067 80 101097 0 FreeSans 240 0 0 0 B[3]
port 11 nsew signal input
flabel metal3 s 0 100251 80 100281 0 FreeSans 240 0 0 0 B[4]
port 12 nsew signal input
flabel metal3 s 0 99571 80 99601 0 FreeSans 240 0 0 0 B[5]
port 13 nsew signal input
flabel metal3 s 0 99299 80 99329 0 FreeSans 240 0 0 0 B[6]
port 14 nsew signal input
flabel metal3 s 0 101475 80 101505 0 FreeSans 240 0 0 0 B[7]
port 15 nsew signal input
flabel metal3 s 0 100387 80 100417 0 FreeSans 240 0 0 0 Cin
port 16 nsew signal input
flabel metal3 s 0 99435 80 99465 0 FreeSans 240 0 0 0 Cout
port 17 nsew signal output
flabel metal4 s 215 0 245 80 0 FreeSans 240 90 0 0 VDD
port 18 nsew signal input
flabel metal4 s 399 0 429 80 0 FreeSans 240 90 0 0 VSS
port 19 nsew signal input
flabel metal3 s 0 98755 80 98785 0 FreeSans 240 0 0 0 Y[0]
port 20 nsew signal output
flabel metal3 s 0 101203 80 101233 0 FreeSans 240 0 0 0 Y[1]
port 21 nsew signal output
flabel metal3 s 0 101611 80 101641 0 FreeSans 240 0 0 0 Y[2]
port 22 nsew signal output
flabel metal3 s 0 98483 80 98513 0 FreeSans 240 0 0 0 Y[3]
port 23 nsew signal output
flabel metal3 s 0 101339 80 101369 0 FreeSans 240 0 0 0 Y[4]
port 24 nsew signal output
flabel metal3 s 0 100115 80 100145 0 FreeSans 240 0 0 0 Y[5]
port 25 nsew signal output
flabel metal3 s 0 99027 80 99057 0 FreeSans 240 0 0 0 Y[6]
port 26 nsew signal output
flabel metal3 s 0 99163 80 99193 0 FreeSans 240 0 0 0 Y[7]
port 27 nsew signal output
rlabel space 13778 95082 24901 196862 6 help
<< properties >>
string FIXED_BBOX 0 0 200000 200000
<< end >>
