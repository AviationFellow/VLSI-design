******************************************************
* Gate-level SPICE netlist for 8-bit CLA (Sky130)
******************************************************

* Include standard cell library
.include "/home/arumukamganesmoorthe/tools/open_pdks/sky130/sky130A/libs.ref/sky130_fd_sc_hd/spice/sky130_fd_sc_hd.spice"

*-----------------------------------------------------
* Define power supplies
*-----------------------------------------------------
VDD VDD 0 DC 1.8V
VSS VSS 0 DC 0V

*-----------------------------------------------------
* 4-bit CLA Subcircuit
*-----------------------------------------------------
* Node order: A B Cin VDD VSS S0 S1 S2 S3 Cout
.SUBCKT CLA4bit A0 A1 A2 A3 B0 B1 B2 B3 Cin VDD VSS S0 S1 S2 S3 Cout

* Internal carry wires
W0 W1 W2

* XOR/XNOR and majority gates with VDD/VSS connections
X0 B0 A0 VDD VSS W0 sky130_fd_sc_hd__xnor2_1
X1 B0 A0 Cin VDD VSS W1 sky130_fd_sc_hd__maj3_1

X2 B1 A1 VDD VSS W1 W2 sky130_fd_sc_hd__xnor2_1
X3 B1 A1 W1 VDD VSS W2 sky130_fd_sc_hd__maj3_1

X4 B2 A2 VDD VSS W2 W0 sky130_fd_sc_hd__xnor2_1
X5 B2 A2 W2 VDD VSS W0 sky130_fd_sc_hd__maj3_1

X6 B3 A3 VDD VSS W0 W1 sky130_fd_sc_hd__xnor2_1
X7 B3 A3 W0 VDD VSS Cout sky130_fd_sc_hd__maj3_1

* Final sum outputs
X8 Cin W0 VDD VSS S0 sky130_fd_sc_hd__xnor2_1
X9 W1 W2 VDD VSS S1 sky130_fd_sc_hd__xnor2_1
X10 W2 W0 VDD VSS S2 sky130_fd_sc_hd__xnor2_1
X11 W1 W1 VDD VSS S3 sky130_fd_sc_hd__xnor2_1

.ENDS CLA4bit

*-----------------------------------------------------
* 8-bit Adder Subcircuit
*-----------------------------------------------------
* Node order: A0..A7 B0..B7 Cin VDD VSS Y0..Y7 Cout
.SUBCKT eb_adder A0 A1 A2 A3 A4 A5 A6 A7 B0 B1 B2 B3 B4 B5 B6 B7 Cin VDD VSS \
                 Y0 Y1 Y2 Y3 Y4 Y5 Y6 Y7 Cout

* Internal carry between lower and upper 4-bit CLA
WIRE x

XLOW  A0 A1 A2 A3 B0 B1 B2 B3 Cin VDD VSS Y0 Y1 Y2 Y3 x CLA4bit
XUPP  A4 A5 A6 A7 B4 B5 B6 B7 x VDD VSS Y4 Y5 Y6 Y7 Cout CLA4bit

.ENDS eb_adder

*-----------------------------------------------------
* Top-level instantiation
*-----------------------------------------------------
* Inputs
VIN_A0 A0 0 DC 0
VIN_A1 A1 0 DC 0
VIN_A2 A2 0 DC 0
VIN_A3 A3 0 DC 0
VIN_A4 A4 0 DC 0
VIN_A5 A5 0 DC 0
VIN_A6 A6 0 DC 0
VIN_A7 A7 0 DC 0

VIN_B0 B0 0 DC 0
VIN_B1 B1 0 DC 0
VIN_B2 B2 0 DC 0
VIN_B3 B3 0 DC 0
VIN_B4 B4 0 DC 0
VIN_B5 B5 0 DC 0
VIN_B6 B6 0 DC 0
VIN_B7 B7 0 DC 0

VIN_Cin Cin 0 DC 0

* Instantiate the 8-bit adder
XCLA A0 A1 A2 A3 A4 A5 A6 A7 \
      B0 B1 B2 B3 B4 B5 B6 B7 \
      Cin VDD VSS \
      Y0 Y1 Y2 Y3 Y4 Y5 Y6 Y7 Cout \
      eb_adder

*-----------------------------------------------------
* Simulation commands
*-----------------------------------------------------
* Define outputs to monitor
.control
  * Print all outputs
  print V(Y0) V(Y1) V(Y2) V(Y3) V(Y4) V(Y5) V(Y6) V(Y7) V(Cout)
  * Run a DC operating point analysis
  op
  * End control block
.endc

.end

