module vedic1 (a,
    b,
    c);
 input [15:0] a;
 input [15:0] b;
 output [31:0] c;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire \lastadder/Cout ;
 wire \lastadder/ksa32/_000_ ;
 wire \lastadder/ksa32/_001_ ;
 wire \lastadder/ksa32/_002_ ;
 wire \lastadder/ksa32/_003_ ;
 wire \lastadder/ksa32/_004_ ;
 wire \lastadder/ksa32/_005_ ;
 wire \lastadder/ksa32/_006_ ;
 wire \lastadder/ksa32/_007_ ;
 wire \lastadder/ksa32/_008_ ;
 wire \lastadder/ksa32/_009_ ;
 wire \lastadder/ksa32/_010_ ;
 wire \lastadder/ksa32/_011_ ;
 wire \lastadder/ksa32/_012_ ;
 wire \lastadder/ksa32/_013_ ;
 wire \lastadder/ksa32/_014_ ;
 wire \lastadder/ksa32/_015_ ;
 wire \lastadder/ksa32/_016_ ;
 wire \lastadder/ksa32/_017_ ;
 wire \lastadder/ksa32/_018_ ;
 wire \lastadder/ksa32/_019_ ;
 wire \lastadder/ksa32/_020_ ;
 wire \lastadder/ksa32/_021_ ;
 wire \lastadder/ksa32/_022_ ;
 wire \lastadder/ksa32/_023_ ;
 wire \lastadder/ksa32/_024_ ;
 wire \lastadder/ksa32/_025_ ;
 wire \lastadder/ksa32/_026_ ;
 wire \lastadder/ksa32/_027_ ;
 wire \lastadder/ksa32/_028_ ;
 wire \lastadder/ksa32/_029_ ;
 wire \lastadder/ksa32/_030_ ;
 wire \lastadder/ksa32/_031_ ;
 wire \lastadder/ksa32/_032_ ;
 wire \lastadder/ksa32/_033_ ;
 wire \lastadder/ksa32/_034_ ;
 wire \lastadder/ksa32/_035_ ;
 wire \lastadder/ksa32/_036_ ;
 wire \lastadder/ksa32/_037_ ;
 wire \lastadder/ksa32/_038_ ;
 wire \lastadder/ksa32/_039_ ;
 wire \lastadder/ksa32/_040_ ;
 wire \lastadder/ksa32/_041_ ;
 wire \lastadder/ksa32/_042_ ;
 wire \lastadder/ksa32/_043_ ;
 wire \lastadder/ksa32/_044_ ;
 wire \lastadder/ksa32/_045_ ;
 wire \lastadder/ksa32/_046_ ;
 wire \lastadder/ksa32/_047_ ;
 wire \lastadder/ksa32/_048_ ;
 wire \lastadder/ksa32/_049_ ;
 wire \lastadder/ksa32/_050_ ;
 wire \lastadder/ksa32/_051_ ;
 wire \lastadder/ksa32/_052_ ;
 wire \lastadder/ksa32/_053_ ;
 wire \lastadder/ksa32/_054_ ;
 wire \lastadder/ksa32/_055_ ;
 wire \lastadder/ksa32/_056_ ;
 wire \lastadder/ksa32/_057_ ;
 wire \lastadder/ksa32/_058_ ;
 wire \lastadder/ksa32/_059_ ;
 wire \lastadder/ksa32/_060_ ;
 wire \lastadder/ksa32/_061_ ;
 wire \lastadder/ksa32/_062_ ;
 wire \lastadder/ksa32/_063_ ;
 wire \lastadder/ksa32/_064_ ;
 wire \lastadder/ksa32/_065_ ;
 wire \lastadder/ksa32/_066_ ;
 wire \lastadder/ksa32/_067_ ;
 wire \lastadder/ksa32/_068_ ;
 wire \lastadder/ksa32/_069_ ;
 wire \lastadder/ksa32/_070_ ;
 wire \lastadder/ksa32/_071_ ;
 wire \lastadder/ksa32/_072_ ;
 wire \lastadder/ksa32/_073_ ;
 wire \lastadder/ksa32/_074_ ;
 wire \lastadder/ksa32/_075_ ;
 wire \lastadder/ksa32/_076_ ;
 wire \lastadder/ksa32/_077_ ;
 wire \lastadder/ksa32/_078_ ;
 wire \lastadder/ksa32/_079_ ;
 wire \lastadder/ksa32/_080_ ;
 wire \lastadder/ksa32/_081_ ;
 wire \lastadder/ksa32/_082_ ;
 wire \lastadder/ksa32/_083_ ;
 wire \lastadder/ksa32/_084_ ;
 wire \lastadder/ksa32/_085_ ;
 wire \lastadder/ksa32/_086_ ;
 wire \lastadder/ksa32/_087_ ;
 wire \lastadder/ksa32/_088_ ;
 wire \lastadder/ksa32/_089_ ;
 wire \lastadder/ksa32/_090_ ;
 wire \lastadder/ksa32/_091_ ;
 wire \lastadder/ksa32/_092_ ;
 wire \lastadder/ksa32/_093_ ;
 wire \lastadder/ksa32/_094_ ;
 wire \lastadder/ksa32/_095_ ;
 wire \lastadder/ksa32/_096_ ;
 wire \lastadder/ksa32/_097_ ;
 wire \lastadder/ksa32/_098_ ;
 wire \lastadder/ksa32/_099_ ;
 wire \lastadder/ksa32/_100_ ;
 wire \lastadder/ksa32/_101_ ;
 wire \lastadder/ksa32/_102_ ;
 wire \lastadder/ksa32/_103_ ;
 wire \lastadder/ksa32/_104_ ;
 wire \lastadder/ksa32/_105_ ;
 wire \lastadder/ksa32/_106_ ;
 wire \lastadder/ksa32/_107_ ;
 wire \lastadder/ksa32/_108_ ;
 wire \lastadder/ksa32/_109_ ;
 wire \lastadder/ksa32/_110_ ;
 wire \lastadder/ksa32/_111_ ;
 wire \lastadder/ksa32/_112_ ;
 wire \lastadder/ksa32/_113_ ;
 wire \lastadder/ksa32/_114_ ;
 wire \lastadder/ksa32/_115_ ;
 wire \lastadder/ksa32/_116_ ;
 wire \lastadder/ksa32/_117_ ;
 wire \lastadder/ksa32/_118_ ;
 wire \lastadder/ksa32/_119_ ;
 wire \lastadder/ksa32/_120_ ;
 wire \lastadder/ksa32/_121_ ;
 wire \lastadder/ksa32/_122_ ;
 wire \lastadder/ksa32/_123_ ;
 wire \lastadder/ksa32/_124_ ;
 wire \lastadder/ksa32/_125_ ;
 wire \lastadder/ksa32/_126_ ;
 wire \lastadder/ksa32/_127_ ;
 wire \lastadder/ksa32/_128_ ;
 wire \lastadder/ksa32/_129_ ;
 wire \lastadder/ksa32/_130_ ;
 wire \lastadder/ksa32/_131_ ;
 wire \lastadder/ksa32/_132_ ;
 wire \lastadder/ksa32/_133_ ;
 wire \lastadder/ksa32/_134_ ;
 wire \lastadder/ksa32/_135_ ;
 wire \lastadder/ksa32/_136_ ;
 wire \lastadder/ksa32/_137_ ;
 wire \lastadder/ksa32/_138_ ;
 wire \lastadder/ksa32/_139_ ;
 wire \lastadder/ksa32/_140_ ;
 wire \lastadder/ksa32/_141_ ;
 wire \lastadder/ksa32/_142_ ;
 wire \lastadder/ksa32/_143_ ;
 wire \lastadder/ksa32/_144_ ;
 wire \lastadder/ksa32/_145_ ;
 wire \lastadder/ksa32/_146_ ;
 wire \lastadder/ksa32/_147_ ;
 wire \lastadder/ksa32/_148_ ;
 wire \lastadder/ksa32/_149_ ;
 wire \lastadder/ksa32/_150_ ;
 wire \lastadder/ksa32/_151_ ;
 wire \lastadder/ksa32/_152_ ;
 wire \lastadder/ksa32/_153_ ;
 wire \lastadder/ksa32/_154_ ;
 wire \lastadder/ksa32/_155_ ;
 wire \lastadder/ksa32/_156_ ;
 wire \lastadder/ksa32/_157_ ;
 wire \lastadder/ksa32/_158_ ;
 wire \lastadder/ksa32/_159_ ;
 wire \lastadder/ksa32/_160_ ;
 wire \lastadder/ksa32/_161_ ;
 wire \lastadder/ksa32/_162_ ;
 wire sign;
 wire \v0/_00_ ;
 wire \v0/_01_ ;
 wire \v0/_02_ ;
 wire \v0/_03_ ;
 wire \v0/_04_ ;
 wire \v0/_05_ ;
 wire \v0/_06_ ;
 wire \v0/_07_ ;
 wire \v0/_08_ ;
 wire \v0/_09_ ;
 wire \v0/_10_ ;
 wire \v0/_11_ ;
 wire \v0/_12_ ;
 wire \v0/_13_ ;
 wire \v0/_14_ ;
 wire \v0/_15_ ;
 wire \v0/_16_ ;
 wire \v0/_17_ ;
 wire \v0/_18_ ;
 wire \v0/_19_ ;
 wire \v0/_20_ ;
 wire \v0/_21_ ;
 wire \v0/_22_ ;
 wire \v0/_23_ ;
 wire \v0/_24_ ;
 wire \v0/_25_ ;
 wire \v0/_26_ ;
 wire \v0/_27_ ;
 wire \v0/_28_ ;
 wire \v0/_29_ ;
 wire \v0/_30_ ;
 wire \v0/_31_ ;
 wire \v0/_32_ ;
 wire \v0/_33_ ;
 wire \v0/_34_ ;
 wire \v0/z1/_00_ ;
 wire \v0/z1/_01_ ;
 wire \v0/z1/_02_ ;
 wire \v0/z1/_03_ ;
 wire \v0/z1/_04_ ;
 wire \v0/z1/_05_ ;
 wire \v0/z1/_06_ ;
 wire \v0/z1/_07_ ;
 wire \v0/z1/_08_ ;
 wire \v0/z1/_09_ ;
 wire \v0/z1/_10_ ;
 wire \v0/z1/_11_ ;
 wire \v0/z1/_12_ ;
 wire \v0/z1/_13_ ;
 wire \v0/z1/_14_ ;
 wire \v0/z1/_15_ ;
 wire \v0/z1/_16_ ;
 wire \v0/z1/_17_ ;
 wire \v0/z1/_18_ ;
 wire \v0/z1/z1/_00_ ;
 wire \v0/z1/z1/_01_ ;
 wire \v0/z1/z1/_02_ ;
 wire \v0/z1/z1/_03_ ;
 wire \v0/z1/z1/_04_ ;
 wire \v0/z1/z1/_05_ ;
 wire \v0/z1/z1/_06_ ;
 wire \v0/z1/z1/_07_ ;
 wire \v0/z1/z1/_08_ ;
 wire \v0/z1/z1/_09_ ;
 wire \v0/z1/z1/_10_ ;
 wire \v0/z1/z1/z5/Cout ;
 wire \v0/z1/z1/z5/_00_ ;
 wire \v0/z1/z1/z5/_01_ ;
 wire \v0/z1/z1/z5/_02_ ;
 wire \v0/z1/z1/z5/_03_ ;
 wire \v0/z1/z1/z5/_04_ ;
 wire \v0/z1/z1/z5/_05_ ;
 wire \v0/z1/z1/z5/_06_ ;
 wire \v0/z1/z1/z6/Cout ;
 wire \v0/z1/z1/z6/_00_ ;
 wire \v0/z1/z1/z6/_01_ ;
 wire \v0/z1/z1/z6/_02_ ;
 wire \v0/z1/z1/z6/_03_ ;
 wire \v0/z1/z1/z6/_04_ ;
 wire \v0/z1/z1/z6/_05_ ;
 wire \v0/z1/z1/z6/_06_ ;
 wire \v0/z1/z1/z6/_07_ ;
 wire \v0/z1/z1/z6/_08_ ;
 wire \v0/z1/z1/z6/_09_ ;
 wire \v0/z1/z1/z6/_10_ ;
 wire \v0/z1/z1/z6/_11_ ;
 wire \v0/z1/z1/z6/_12_ ;
 wire \v0/z1/z1/z6/_13_ ;
 wire \v0/z1/z1/z6/_14_ ;
 wire \v0/z1/z1/z6/_15_ ;
 wire \v0/z1/z1/z6/_16_ ;
 wire \v0/z1/z1/z6/_17_ ;
 wire \v0/z1/z1/z6/_18_ ;
 wire \v0/z1/z1/z7/Cout ;
 wire \v0/z1/z1/z7/_00_ ;
 wire \v0/z1/z1/z7/_01_ ;
 wire \v0/z1/z1/z7/_02_ ;
 wire \v0/z1/z1/z7/_03_ ;
 wire \v0/z1/z1/z7/_04_ ;
 wire \v0/z1/z1/z7/_05_ ;
 wire \v0/z1/z1/z7/_06_ ;
 wire \v0/z1/z1/z7/_07_ ;
 wire \v0/z1/z1/z7/_08_ ;
 wire \v0/z1/z1/z7/_09_ ;
 wire \v0/z1/z1/z7/_10_ ;
 wire \v0/z1/z1/z7/_11_ ;
 wire \v0/z1/z1/z7/_12_ ;
 wire \v0/z1/z1/z7/_13_ ;
 wire \v0/z1/z1/z7/_14_ ;
 wire \v0/z1/z1/z7/_15_ ;
 wire \v0/z1/z1/z7/_16_ ;
 wire \v0/z1/z1/z7/_17_ ;
 wire \v0/z1/z1/z7/_18_ ;
 wire \v0/z1/z2/_00_ ;
 wire \v0/z1/z2/_01_ ;
 wire \v0/z1/z2/_02_ ;
 wire \v0/z1/z2/_03_ ;
 wire \v0/z1/z2/_04_ ;
 wire \v0/z1/z2/_05_ ;
 wire \v0/z1/z2/_06_ ;
 wire \v0/z1/z2/_07_ ;
 wire \v0/z1/z2/_08_ ;
 wire \v0/z1/z2/_09_ ;
 wire \v0/z1/z2/_10_ ;
 wire \v0/z1/z2/z5/Cout ;
 wire \v0/z1/z2/z5/_00_ ;
 wire \v0/z1/z2/z5/_01_ ;
 wire \v0/z1/z2/z5/_02_ ;
 wire \v0/z1/z2/z5/_03_ ;
 wire \v0/z1/z2/z5/_04_ ;
 wire \v0/z1/z2/z5/_05_ ;
 wire \v0/z1/z2/z5/_06_ ;
 wire \v0/z1/z2/z6/Cout ;
 wire \v0/z1/z2/z6/_00_ ;
 wire \v0/z1/z2/z6/_01_ ;
 wire \v0/z1/z2/z6/_02_ ;
 wire \v0/z1/z2/z6/_03_ ;
 wire \v0/z1/z2/z6/_04_ ;
 wire \v0/z1/z2/z6/_05_ ;
 wire \v0/z1/z2/z6/_06_ ;
 wire \v0/z1/z2/z6/_07_ ;
 wire \v0/z1/z2/z6/_08_ ;
 wire \v0/z1/z2/z6/_09_ ;
 wire \v0/z1/z2/z6/_10_ ;
 wire \v0/z1/z2/z6/_11_ ;
 wire \v0/z1/z2/z6/_12_ ;
 wire \v0/z1/z2/z6/_13_ ;
 wire \v0/z1/z2/z6/_14_ ;
 wire \v0/z1/z2/z6/_15_ ;
 wire \v0/z1/z2/z6/_16_ ;
 wire \v0/z1/z2/z6/_17_ ;
 wire \v0/z1/z2/z6/_18_ ;
 wire \v0/z1/z2/z7/Cout ;
 wire \v0/z1/z2/z7/_00_ ;
 wire \v0/z1/z2/z7/_01_ ;
 wire \v0/z1/z2/z7/_02_ ;
 wire \v0/z1/z2/z7/_03_ ;
 wire \v0/z1/z2/z7/_04_ ;
 wire \v0/z1/z2/z7/_05_ ;
 wire \v0/z1/z2/z7/_06_ ;
 wire \v0/z1/z2/z7/_07_ ;
 wire \v0/z1/z2/z7/_08_ ;
 wire \v0/z1/z2/z7/_09_ ;
 wire \v0/z1/z2/z7/_10_ ;
 wire \v0/z1/z2/z7/_11_ ;
 wire \v0/z1/z2/z7/_12_ ;
 wire \v0/z1/z2/z7/_13_ ;
 wire \v0/z1/z2/z7/_14_ ;
 wire \v0/z1/z2/z7/_15_ ;
 wire \v0/z1/z2/z7/_16_ ;
 wire \v0/z1/z2/z7/_17_ ;
 wire \v0/z1/z2/z7/_18_ ;
 wire \v0/z1/z3/_00_ ;
 wire \v0/z1/z3/_01_ ;
 wire \v0/z1/z3/_02_ ;
 wire \v0/z1/z3/_03_ ;
 wire \v0/z1/z3/_04_ ;
 wire \v0/z1/z3/_05_ ;
 wire \v0/z1/z3/_06_ ;
 wire \v0/z1/z3/_07_ ;
 wire \v0/z1/z3/_08_ ;
 wire \v0/z1/z3/_09_ ;
 wire \v0/z1/z3/_10_ ;
 wire \v0/z1/z3/z5/Cout ;
 wire \v0/z1/z3/z5/_00_ ;
 wire \v0/z1/z3/z5/_01_ ;
 wire \v0/z1/z3/z5/_02_ ;
 wire \v0/z1/z3/z5/_03_ ;
 wire \v0/z1/z3/z5/_04_ ;
 wire \v0/z1/z3/z5/_05_ ;
 wire \v0/z1/z3/z5/_06_ ;
 wire \v0/z1/z3/z6/Cout ;
 wire \v0/z1/z3/z6/_00_ ;
 wire \v0/z1/z3/z6/_01_ ;
 wire \v0/z1/z3/z6/_02_ ;
 wire \v0/z1/z3/z6/_03_ ;
 wire \v0/z1/z3/z6/_04_ ;
 wire \v0/z1/z3/z6/_05_ ;
 wire \v0/z1/z3/z6/_06_ ;
 wire \v0/z1/z3/z6/_07_ ;
 wire \v0/z1/z3/z6/_08_ ;
 wire \v0/z1/z3/z6/_09_ ;
 wire \v0/z1/z3/z6/_10_ ;
 wire \v0/z1/z3/z6/_11_ ;
 wire \v0/z1/z3/z6/_12_ ;
 wire \v0/z1/z3/z6/_13_ ;
 wire \v0/z1/z3/z6/_14_ ;
 wire \v0/z1/z3/z6/_15_ ;
 wire \v0/z1/z3/z6/_16_ ;
 wire \v0/z1/z3/z6/_17_ ;
 wire \v0/z1/z3/z6/_18_ ;
 wire \v0/z1/z3/z7/Cout ;
 wire \v0/z1/z3/z7/_00_ ;
 wire \v0/z1/z3/z7/_01_ ;
 wire \v0/z1/z3/z7/_02_ ;
 wire \v0/z1/z3/z7/_03_ ;
 wire \v0/z1/z3/z7/_04_ ;
 wire \v0/z1/z3/z7/_05_ ;
 wire \v0/z1/z3/z7/_06_ ;
 wire \v0/z1/z3/z7/_07_ ;
 wire \v0/z1/z3/z7/_08_ ;
 wire \v0/z1/z3/z7/_09_ ;
 wire \v0/z1/z3/z7/_10_ ;
 wire \v0/z1/z3/z7/_11_ ;
 wire \v0/z1/z3/z7/_12_ ;
 wire \v0/z1/z3/z7/_13_ ;
 wire \v0/z1/z3/z7/_14_ ;
 wire \v0/z1/z3/z7/_15_ ;
 wire \v0/z1/z3/z7/_16_ ;
 wire \v0/z1/z3/z7/_17_ ;
 wire \v0/z1/z3/z7/_18_ ;
 wire \v0/z1/z4/_00_ ;
 wire \v0/z1/z4/_01_ ;
 wire \v0/z1/z4/_02_ ;
 wire \v0/z1/z4/_03_ ;
 wire \v0/z1/z4/_04_ ;
 wire \v0/z1/z4/_05_ ;
 wire \v0/z1/z4/_06_ ;
 wire \v0/z1/z4/_07_ ;
 wire \v0/z1/z4/_08_ ;
 wire \v0/z1/z4/_09_ ;
 wire \v0/z1/z4/_10_ ;
 wire \v0/z1/z4/z5/Cout ;
 wire \v0/z1/z4/z5/_00_ ;
 wire \v0/z1/z4/z5/_01_ ;
 wire \v0/z1/z4/z5/_02_ ;
 wire \v0/z1/z4/z5/_03_ ;
 wire \v0/z1/z4/z5/_04_ ;
 wire \v0/z1/z4/z5/_05_ ;
 wire \v0/z1/z4/z5/_06_ ;
 wire \v0/z1/z4/z6/Cout ;
 wire \v0/z1/z4/z6/_00_ ;
 wire \v0/z1/z4/z6/_01_ ;
 wire \v0/z1/z4/z6/_02_ ;
 wire \v0/z1/z4/z6/_03_ ;
 wire \v0/z1/z4/z6/_04_ ;
 wire \v0/z1/z4/z6/_05_ ;
 wire \v0/z1/z4/z6/_06_ ;
 wire \v0/z1/z4/z6/_07_ ;
 wire \v0/z1/z4/z6/_08_ ;
 wire \v0/z1/z4/z6/_09_ ;
 wire \v0/z1/z4/z6/_10_ ;
 wire \v0/z1/z4/z6/_11_ ;
 wire \v0/z1/z4/z6/_12_ ;
 wire \v0/z1/z4/z6/_13_ ;
 wire \v0/z1/z4/z6/_14_ ;
 wire \v0/z1/z4/z6/_15_ ;
 wire \v0/z1/z4/z6/_16_ ;
 wire \v0/z1/z4/z6/_17_ ;
 wire \v0/z1/z4/z6/_18_ ;
 wire \v0/z1/z4/z7/Cout ;
 wire \v0/z1/z4/z7/_00_ ;
 wire \v0/z1/z4/z7/_01_ ;
 wire \v0/z1/z4/z7/_02_ ;
 wire \v0/z1/z4/z7/_03_ ;
 wire \v0/z1/z4/z7/_04_ ;
 wire \v0/z1/z4/z7/_05_ ;
 wire \v0/z1/z4/z7/_06_ ;
 wire \v0/z1/z4/z7/_07_ ;
 wire \v0/z1/z4/z7/_08_ ;
 wire \v0/z1/z4/z7/_09_ ;
 wire \v0/z1/z4/z7/_10_ ;
 wire \v0/z1/z4/z7/_11_ ;
 wire \v0/z1/z4/z7/_12_ ;
 wire \v0/z1/z4/z7/_13_ ;
 wire \v0/z1/z4/z7/_14_ ;
 wire \v0/z1/z4/z7/_15_ ;
 wire \v0/z1/z4/z7/_16_ ;
 wire \v0/z1/z4/z7/_17_ ;
 wire \v0/z1/z4/z7/_18_ ;
 wire \v0/z1/z5/Cout ;
 wire \v0/z1/z5/_00_ ;
 wire \v0/z1/z5/_01_ ;
 wire \v0/z1/z5/_02_ ;
 wire \v0/z1/z5/_03_ ;
 wire \v0/z1/z5/_04_ ;
 wire \v0/z1/z5/_05_ ;
 wire \v0/z1/z5/_06_ ;
 wire \v0/z1/z5/_07_ ;
 wire \v0/z1/z5/_08_ ;
 wire \v0/z1/z5/_09_ ;
 wire \v0/z1/z5/_10_ ;
 wire \v0/z1/z5/_11_ ;
 wire \v0/z1/z5/_12_ ;
 wire \v0/z1/z5/_13_ ;
 wire \v0/z1/z5/_14_ ;
 wire \v0/z1/z5/_15_ ;
 wire \v0/z1/z5/_16_ ;
 wire \v0/z1/z5/_17_ ;
 wire \v0/z1/z5/_18_ ;
 wire \v0/z1/z5/_19_ ;
 wire \v0/z1/z5/_20_ ;
 wire \v0/z1/z5/_21_ ;
 wire \v0/z1/z5/_22_ ;
 wire \v0/z1/z5/_23_ ;
 wire \v0/z1/z5/_24_ ;
 wire \v0/z1/z5/_25_ ;
 wire \v0/z1/z5/_26_ ;
 wire \v0/z1/z6/Cout ;
 wire \v0/z1/z6/_000_ ;
 wire \v0/z1/z6/_001_ ;
 wire \v0/z1/z6/_002_ ;
 wire \v0/z1/z6/_003_ ;
 wire \v0/z1/z6/_004_ ;
 wire \v0/z1/z6/_005_ ;
 wire \v0/z1/z6/_006_ ;
 wire \v0/z1/z6/_007_ ;
 wire \v0/z1/z6/_008_ ;
 wire \v0/z1/z6/_009_ ;
 wire \v0/z1/z6/_010_ ;
 wire \v0/z1/z6/_011_ ;
 wire \v0/z1/z6/_012_ ;
 wire \v0/z1/z6/_013_ ;
 wire \v0/z1/z6/_014_ ;
 wire \v0/z1/z6/_015_ ;
 wire \v0/z1/z6/_016_ ;
 wire \v0/z1/z6/_017_ ;
 wire \v0/z1/z6/_018_ ;
 wire \v0/z1/z6/_019_ ;
 wire \v0/z1/z6/_020_ ;
 wire \v0/z1/z6/_021_ ;
 wire \v0/z1/z6/_022_ ;
 wire \v0/z1/z6/_023_ ;
 wire \v0/z1/z6/_024_ ;
 wire \v0/z1/z6/_025_ ;
 wire \v0/z1/z6/_026_ ;
 wire \v0/z1/z6/_027_ ;
 wire \v0/z1/z6/_028_ ;
 wire \v0/z1/z6/_029_ ;
 wire \v0/z1/z6/_030_ ;
 wire \v0/z1/z6/_031_ ;
 wire \v0/z1/z6/_032_ ;
 wire \v0/z1/z6/_033_ ;
 wire \v0/z1/z6/_034_ ;
 wire \v0/z1/z6/_035_ ;
 wire \v0/z1/z6/_036_ ;
 wire \v0/z1/z6/_037_ ;
 wire \v0/z1/z6/_038_ ;
 wire \v0/z1/z6/_039_ ;
 wire \v0/z1/z6/_040_ ;
 wire \v0/z1/z6/_041_ ;
 wire \v0/z1/z6/_042_ ;
 wire \v0/z1/z6/_043_ ;
 wire \v0/z1/z6/_044_ ;
 wire \v0/z1/z6/_045_ ;
 wire \v0/z1/z6/_046_ ;
 wire \v0/z1/z6/_047_ ;
 wire \v0/z1/z6/_048_ ;
 wire \v0/z1/z6/_049_ ;
 wire \v0/z1/z7/Cout ;
 wire \v0/z1/z7/_000_ ;
 wire \v0/z1/z7/_001_ ;
 wire \v0/z1/z7/_002_ ;
 wire \v0/z1/z7/_003_ ;
 wire \v0/z1/z7/_004_ ;
 wire \v0/z1/z7/_005_ ;
 wire \v0/z1/z7/_006_ ;
 wire \v0/z1/z7/_007_ ;
 wire \v0/z1/z7/_008_ ;
 wire \v0/z1/z7/_009_ ;
 wire \v0/z1/z7/_010_ ;
 wire \v0/z1/z7/_011_ ;
 wire \v0/z1/z7/_012_ ;
 wire \v0/z1/z7/_013_ ;
 wire \v0/z1/z7/_014_ ;
 wire \v0/z1/z7/_015_ ;
 wire \v0/z1/z7/_016_ ;
 wire \v0/z1/z7/_017_ ;
 wire \v0/z1/z7/_018_ ;
 wire \v0/z1/z7/_019_ ;
 wire \v0/z1/z7/_020_ ;
 wire \v0/z1/z7/_021_ ;
 wire \v0/z1/z7/_022_ ;
 wire \v0/z1/z7/_023_ ;
 wire \v0/z1/z7/_024_ ;
 wire \v0/z1/z7/_025_ ;
 wire \v0/z1/z7/_026_ ;
 wire \v0/z1/z7/_027_ ;
 wire \v0/z1/z7/_028_ ;
 wire \v0/z1/z7/_029_ ;
 wire \v0/z1/z7/_030_ ;
 wire \v0/z1/z7/_031_ ;
 wire \v0/z1/z7/_032_ ;
 wire \v0/z1/z7/_033_ ;
 wire \v0/z1/z7/_034_ ;
 wire \v0/z1/z7/_035_ ;
 wire \v0/z1/z7/_036_ ;
 wire \v0/z1/z7/_037_ ;
 wire \v0/z1/z7/_038_ ;
 wire \v0/z1/z7/_039_ ;
 wire \v0/z1/z7/_040_ ;
 wire \v0/z1/z7/_041_ ;
 wire \v0/z1/z7/_042_ ;
 wire \v0/z1/z7/_043_ ;
 wire \v0/z1/z7/_044_ ;
 wire \v0/z1/z7/_045_ ;
 wire \v0/z1/z7/_046_ ;
 wire \v0/z1/z7/_047_ ;
 wire \v0/z1/z7/_048_ ;
 wire \v0/z1/z7/_049_ ;
 wire \v0/z2/_00_ ;
 wire \v0/z2/_01_ ;
 wire \v0/z2/_02_ ;
 wire \v0/z2/_03_ ;
 wire \v0/z2/_04_ ;
 wire \v0/z2/_05_ ;
 wire \v0/z2/_06_ ;
 wire \v0/z2/_07_ ;
 wire \v0/z2/_08_ ;
 wire \v0/z2/_09_ ;
 wire \v0/z2/_10_ ;
 wire \v0/z2/_11_ ;
 wire \v0/z2/_12_ ;
 wire \v0/z2/_13_ ;
 wire \v0/z2/_14_ ;
 wire \v0/z2/_15_ ;
 wire \v0/z2/_16_ ;
 wire \v0/z2/_17_ ;
 wire \v0/z2/_18_ ;
 wire \v0/z2/z1/_00_ ;
 wire \v0/z2/z1/_01_ ;
 wire \v0/z2/z1/_02_ ;
 wire \v0/z2/z1/_03_ ;
 wire \v0/z2/z1/_04_ ;
 wire \v0/z2/z1/_05_ ;
 wire \v0/z2/z1/_06_ ;
 wire \v0/z2/z1/_07_ ;
 wire \v0/z2/z1/_08_ ;
 wire \v0/z2/z1/_09_ ;
 wire \v0/z2/z1/_10_ ;
 wire \v0/z2/z1/z5/Cout ;
 wire \v0/z2/z1/z5/_00_ ;
 wire \v0/z2/z1/z5/_01_ ;
 wire \v0/z2/z1/z5/_02_ ;
 wire \v0/z2/z1/z5/_03_ ;
 wire \v0/z2/z1/z5/_04_ ;
 wire \v0/z2/z1/z5/_05_ ;
 wire \v0/z2/z1/z5/_06_ ;
 wire \v0/z2/z1/z6/Cout ;
 wire \v0/z2/z1/z6/_00_ ;
 wire \v0/z2/z1/z6/_01_ ;
 wire \v0/z2/z1/z6/_02_ ;
 wire \v0/z2/z1/z6/_03_ ;
 wire \v0/z2/z1/z6/_04_ ;
 wire \v0/z2/z1/z6/_05_ ;
 wire \v0/z2/z1/z6/_06_ ;
 wire \v0/z2/z1/z6/_07_ ;
 wire \v0/z2/z1/z6/_08_ ;
 wire \v0/z2/z1/z6/_09_ ;
 wire \v0/z2/z1/z6/_10_ ;
 wire \v0/z2/z1/z6/_11_ ;
 wire \v0/z2/z1/z6/_12_ ;
 wire \v0/z2/z1/z6/_13_ ;
 wire \v0/z2/z1/z6/_14_ ;
 wire \v0/z2/z1/z6/_15_ ;
 wire \v0/z2/z1/z6/_16_ ;
 wire \v0/z2/z1/z6/_17_ ;
 wire \v0/z2/z1/z6/_18_ ;
 wire \v0/z2/z1/z7/Cout ;
 wire \v0/z2/z1/z7/_00_ ;
 wire \v0/z2/z1/z7/_01_ ;
 wire \v0/z2/z1/z7/_02_ ;
 wire \v0/z2/z1/z7/_03_ ;
 wire \v0/z2/z1/z7/_04_ ;
 wire \v0/z2/z1/z7/_05_ ;
 wire \v0/z2/z1/z7/_06_ ;
 wire \v0/z2/z1/z7/_07_ ;
 wire \v0/z2/z1/z7/_08_ ;
 wire \v0/z2/z1/z7/_09_ ;
 wire \v0/z2/z1/z7/_10_ ;
 wire \v0/z2/z1/z7/_11_ ;
 wire \v0/z2/z1/z7/_12_ ;
 wire \v0/z2/z1/z7/_13_ ;
 wire \v0/z2/z1/z7/_14_ ;
 wire \v0/z2/z1/z7/_15_ ;
 wire \v0/z2/z1/z7/_16_ ;
 wire \v0/z2/z1/z7/_17_ ;
 wire \v0/z2/z1/z7/_18_ ;
 wire \v0/z2/z2/_00_ ;
 wire \v0/z2/z2/_01_ ;
 wire \v0/z2/z2/_02_ ;
 wire \v0/z2/z2/_03_ ;
 wire \v0/z2/z2/_04_ ;
 wire \v0/z2/z2/_05_ ;
 wire \v0/z2/z2/_06_ ;
 wire \v0/z2/z2/_07_ ;
 wire \v0/z2/z2/_08_ ;
 wire \v0/z2/z2/_09_ ;
 wire \v0/z2/z2/_10_ ;
 wire \v0/z2/z2/z5/Cout ;
 wire \v0/z2/z2/z5/_00_ ;
 wire \v0/z2/z2/z5/_01_ ;
 wire \v0/z2/z2/z5/_02_ ;
 wire \v0/z2/z2/z5/_03_ ;
 wire \v0/z2/z2/z5/_04_ ;
 wire \v0/z2/z2/z5/_05_ ;
 wire \v0/z2/z2/z5/_06_ ;
 wire \v0/z2/z2/z6/Cout ;
 wire \v0/z2/z2/z6/_00_ ;
 wire \v0/z2/z2/z6/_01_ ;
 wire \v0/z2/z2/z6/_02_ ;
 wire \v0/z2/z2/z6/_03_ ;
 wire \v0/z2/z2/z6/_04_ ;
 wire \v0/z2/z2/z6/_05_ ;
 wire \v0/z2/z2/z6/_06_ ;
 wire \v0/z2/z2/z6/_07_ ;
 wire \v0/z2/z2/z6/_08_ ;
 wire \v0/z2/z2/z6/_09_ ;
 wire \v0/z2/z2/z6/_10_ ;
 wire \v0/z2/z2/z6/_11_ ;
 wire \v0/z2/z2/z6/_12_ ;
 wire \v0/z2/z2/z6/_13_ ;
 wire \v0/z2/z2/z6/_14_ ;
 wire \v0/z2/z2/z6/_15_ ;
 wire \v0/z2/z2/z6/_16_ ;
 wire \v0/z2/z2/z6/_17_ ;
 wire \v0/z2/z2/z6/_18_ ;
 wire \v0/z2/z2/z7/Cout ;
 wire \v0/z2/z2/z7/_00_ ;
 wire \v0/z2/z2/z7/_01_ ;
 wire \v0/z2/z2/z7/_02_ ;
 wire \v0/z2/z2/z7/_03_ ;
 wire \v0/z2/z2/z7/_04_ ;
 wire \v0/z2/z2/z7/_05_ ;
 wire \v0/z2/z2/z7/_06_ ;
 wire \v0/z2/z2/z7/_07_ ;
 wire \v0/z2/z2/z7/_08_ ;
 wire \v0/z2/z2/z7/_09_ ;
 wire \v0/z2/z2/z7/_10_ ;
 wire \v0/z2/z2/z7/_11_ ;
 wire \v0/z2/z2/z7/_12_ ;
 wire \v0/z2/z2/z7/_13_ ;
 wire \v0/z2/z2/z7/_14_ ;
 wire \v0/z2/z2/z7/_15_ ;
 wire \v0/z2/z2/z7/_16_ ;
 wire \v0/z2/z2/z7/_17_ ;
 wire \v0/z2/z2/z7/_18_ ;
 wire \v0/z2/z3/_00_ ;
 wire \v0/z2/z3/_01_ ;
 wire \v0/z2/z3/_02_ ;
 wire \v0/z2/z3/_03_ ;
 wire \v0/z2/z3/_04_ ;
 wire \v0/z2/z3/_05_ ;
 wire \v0/z2/z3/_06_ ;
 wire \v0/z2/z3/_07_ ;
 wire \v0/z2/z3/_08_ ;
 wire \v0/z2/z3/_09_ ;
 wire \v0/z2/z3/_10_ ;
 wire \v0/z2/z3/z5/Cout ;
 wire \v0/z2/z3/z5/_00_ ;
 wire \v0/z2/z3/z5/_01_ ;
 wire \v0/z2/z3/z5/_02_ ;
 wire \v0/z2/z3/z5/_03_ ;
 wire \v0/z2/z3/z5/_04_ ;
 wire \v0/z2/z3/z5/_05_ ;
 wire \v0/z2/z3/z5/_06_ ;
 wire \v0/z2/z3/z6/Cout ;
 wire \v0/z2/z3/z6/_00_ ;
 wire \v0/z2/z3/z6/_01_ ;
 wire \v0/z2/z3/z6/_02_ ;
 wire \v0/z2/z3/z6/_03_ ;
 wire \v0/z2/z3/z6/_04_ ;
 wire \v0/z2/z3/z6/_05_ ;
 wire \v0/z2/z3/z6/_06_ ;
 wire \v0/z2/z3/z6/_07_ ;
 wire \v0/z2/z3/z6/_08_ ;
 wire \v0/z2/z3/z6/_09_ ;
 wire \v0/z2/z3/z6/_10_ ;
 wire \v0/z2/z3/z6/_11_ ;
 wire \v0/z2/z3/z6/_12_ ;
 wire \v0/z2/z3/z6/_13_ ;
 wire \v0/z2/z3/z6/_14_ ;
 wire \v0/z2/z3/z6/_15_ ;
 wire \v0/z2/z3/z6/_16_ ;
 wire \v0/z2/z3/z6/_17_ ;
 wire \v0/z2/z3/z6/_18_ ;
 wire \v0/z2/z3/z7/Cout ;
 wire \v0/z2/z3/z7/_00_ ;
 wire \v0/z2/z3/z7/_01_ ;
 wire \v0/z2/z3/z7/_02_ ;
 wire \v0/z2/z3/z7/_03_ ;
 wire \v0/z2/z3/z7/_04_ ;
 wire \v0/z2/z3/z7/_05_ ;
 wire \v0/z2/z3/z7/_06_ ;
 wire \v0/z2/z3/z7/_07_ ;
 wire \v0/z2/z3/z7/_08_ ;
 wire \v0/z2/z3/z7/_09_ ;
 wire \v0/z2/z3/z7/_10_ ;
 wire \v0/z2/z3/z7/_11_ ;
 wire \v0/z2/z3/z7/_12_ ;
 wire \v0/z2/z3/z7/_13_ ;
 wire \v0/z2/z3/z7/_14_ ;
 wire \v0/z2/z3/z7/_15_ ;
 wire \v0/z2/z3/z7/_16_ ;
 wire \v0/z2/z3/z7/_17_ ;
 wire \v0/z2/z3/z7/_18_ ;
 wire \v0/z2/z4/_00_ ;
 wire \v0/z2/z4/_01_ ;
 wire \v0/z2/z4/_02_ ;
 wire \v0/z2/z4/_03_ ;
 wire \v0/z2/z4/_04_ ;
 wire \v0/z2/z4/_05_ ;
 wire \v0/z2/z4/_06_ ;
 wire \v0/z2/z4/_07_ ;
 wire \v0/z2/z4/_08_ ;
 wire \v0/z2/z4/_09_ ;
 wire \v0/z2/z4/_10_ ;
 wire \v0/z2/z4/z5/Cout ;
 wire \v0/z2/z4/z5/_00_ ;
 wire \v0/z2/z4/z5/_01_ ;
 wire \v0/z2/z4/z5/_02_ ;
 wire \v0/z2/z4/z5/_03_ ;
 wire \v0/z2/z4/z5/_04_ ;
 wire \v0/z2/z4/z5/_05_ ;
 wire \v0/z2/z4/z5/_06_ ;
 wire \v0/z2/z4/z6/Cout ;
 wire \v0/z2/z4/z6/_00_ ;
 wire \v0/z2/z4/z6/_01_ ;
 wire \v0/z2/z4/z6/_02_ ;
 wire \v0/z2/z4/z6/_03_ ;
 wire \v0/z2/z4/z6/_04_ ;
 wire \v0/z2/z4/z6/_05_ ;
 wire \v0/z2/z4/z6/_06_ ;
 wire \v0/z2/z4/z6/_07_ ;
 wire \v0/z2/z4/z6/_08_ ;
 wire \v0/z2/z4/z6/_09_ ;
 wire \v0/z2/z4/z6/_10_ ;
 wire \v0/z2/z4/z6/_11_ ;
 wire \v0/z2/z4/z6/_12_ ;
 wire \v0/z2/z4/z6/_13_ ;
 wire \v0/z2/z4/z6/_14_ ;
 wire \v0/z2/z4/z6/_15_ ;
 wire \v0/z2/z4/z6/_16_ ;
 wire \v0/z2/z4/z6/_17_ ;
 wire \v0/z2/z4/z6/_18_ ;
 wire \v0/z2/z4/z7/Cout ;
 wire \v0/z2/z4/z7/_00_ ;
 wire \v0/z2/z4/z7/_01_ ;
 wire \v0/z2/z4/z7/_02_ ;
 wire \v0/z2/z4/z7/_03_ ;
 wire \v0/z2/z4/z7/_04_ ;
 wire \v0/z2/z4/z7/_05_ ;
 wire \v0/z2/z4/z7/_06_ ;
 wire \v0/z2/z4/z7/_07_ ;
 wire \v0/z2/z4/z7/_08_ ;
 wire \v0/z2/z4/z7/_09_ ;
 wire \v0/z2/z4/z7/_10_ ;
 wire \v0/z2/z4/z7/_11_ ;
 wire \v0/z2/z4/z7/_12_ ;
 wire \v0/z2/z4/z7/_13_ ;
 wire \v0/z2/z4/z7/_14_ ;
 wire \v0/z2/z4/z7/_15_ ;
 wire \v0/z2/z4/z7/_16_ ;
 wire \v0/z2/z4/z7/_17_ ;
 wire \v0/z2/z4/z7/_18_ ;
 wire \v0/z2/z5/Cout ;
 wire \v0/z2/z5/_00_ ;
 wire \v0/z2/z5/_01_ ;
 wire \v0/z2/z5/_02_ ;
 wire \v0/z2/z5/_03_ ;
 wire \v0/z2/z5/_04_ ;
 wire \v0/z2/z5/_05_ ;
 wire \v0/z2/z5/_06_ ;
 wire \v0/z2/z5/_07_ ;
 wire \v0/z2/z5/_08_ ;
 wire \v0/z2/z5/_09_ ;
 wire \v0/z2/z5/_10_ ;
 wire \v0/z2/z5/_11_ ;
 wire \v0/z2/z5/_12_ ;
 wire \v0/z2/z5/_13_ ;
 wire \v0/z2/z5/_14_ ;
 wire \v0/z2/z5/_15_ ;
 wire \v0/z2/z5/_16_ ;
 wire \v0/z2/z5/_17_ ;
 wire \v0/z2/z5/_18_ ;
 wire \v0/z2/z5/_19_ ;
 wire \v0/z2/z5/_20_ ;
 wire \v0/z2/z5/_21_ ;
 wire \v0/z2/z5/_22_ ;
 wire \v0/z2/z5/_23_ ;
 wire \v0/z2/z5/_24_ ;
 wire \v0/z2/z5/_25_ ;
 wire \v0/z2/z5/_26_ ;
 wire \v0/z2/z6/Cout ;
 wire \v0/z2/z6/_000_ ;
 wire \v0/z2/z6/_001_ ;
 wire \v0/z2/z6/_002_ ;
 wire \v0/z2/z6/_003_ ;
 wire \v0/z2/z6/_004_ ;
 wire \v0/z2/z6/_005_ ;
 wire \v0/z2/z6/_006_ ;
 wire \v0/z2/z6/_007_ ;
 wire \v0/z2/z6/_008_ ;
 wire \v0/z2/z6/_009_ ;
 wire \v0/z2/z6/_010_ ;
 wire \v0/z2/z6/_011_ ;
 wire \v0/z2/z6/_012_ ;
 wire \v0/z2/z6/_013_ ;
 wire \v0/z2/z6/_014_ ;
 wire \v0/z2/z6/_015_ ;
 wire \v0/z2/z6/_016_ ;
 wire \v0/z2/z6/_017_ ;
 wire \v0/z2/z6/_018_ ;
 wire \v0/z2/z6/_019_ ;
 wire \v0/z2/z6/_020_ ;
 wire \v0/z2/z6/_021_ ;
 wire \v0/z2/z6/_022_ ;
 wire \v0/z2/z6/_023_ ;
 wire \v0/z2/z6/_024_ ;
 wire \v0/z2/z6/_025_ ;
 wire \v0/z2/z6/_026_ ;
 wire \v0/z2/z6/_027_ ;
 wire \v0/z2/z6/_028_ ;
 wire \v0/z2/z6/_029_ ;
 wire \v0/z2/z6/_030_ ;
 wire \v0/z2/z6/_031_ ;
 wire \v0/z2/z6/_032_ ;
 wire \v0/z2/z6/_033_ ;
 wire \v0/z2/z6/_034_ ;
 wire \v0/z2/z6/_035_ ;
 wire \v0/z2/z6/_036_ ;
 wire \v0/z2/z6/_037_ ;
 wire \v0/z2/z6/_038_ ;
 wire \v0/z2/z6/_039_ ;
 wire \v0/z2/z6/_040_ ;
 wire \v0/z2/z6/_041_ ;
 wire \v0/z2/z6/_042_ ;
 wire \v0/z2/z6/_043_ ;
 wire \v0/z2/z6/_044_ ;
 wire \v0/z2/z6/_045_ ;
 wire \v0/z2/z6/_046_ ;
 wire \v0/z2/z6/_047_ ;
 wire \v0/z2/z6/_048_ ;
 wire \v0/z2/z6/_049_ ;
 wire \v0/z2/z7/Cout ;
 wire \v0/z2/z7/_000_ ;
 wire \v0/z2/z7/_001_ ;
 wire \v0/z2/z7/_002_ ;
 wire \v0/z2/z7/_003_ ;
 wire \v0/z2/z7/_004_ ;
 wire \v0/z2/z7/_005_ ;
 wire \v0/z2/z7/_006_ ;
 wire \v0/z2/z7/_007_ ;
 wire \v0/z2/z7/_008_ ;
 wire \v0/z2/z7/_009_ ;
 wire \v0/z2/z7/_010_ ;
 wire \v0/z2/z7/_011_ ;
 wire \v0/z2/z7/_012_ ;
 wire \v0/z2/z7/_013_ ;
 wire \v0/z2/z7/_014_ ;
 wire \v0/z2/z7/_015_ ;
 wire \v0/z2/z7/_016_ ;
 wire \v0/z2/z7/_017_ ;
 wire \v0/z2/z7/_018_ ;
 wire \v0/z2/z7/_019_ ;
 wire \v0/z2/z7/_020_ ;
 wire \v0/z2/z7/_021_ ;
 wire \v0/z2/z7/_022_ ;
 wire \v0/z2/z7/_023_ ;
 wire \v0/z2/z7/_024_ ;
 wire \v0/z2/z7/_025_ ;
 wire \v0/z2/z7/_026_ ;
 wire \v0/z2/z7/_027_ ;
 wire \v0/z2/z7/_028_ ;
 wire \v0/z2/z7/_029_ ;
 wire \v0/z2/z7/_030_ ;
 wire \v0/z2/z7/_031_ ;
 wire \v0/z2/z7/_032_ ;
 wire \v0/z2/z7/_033_ ;
 wire \v0/z2/z7/_034_ ;
 wire \v0/z2/z7/_035_ ;
 wire \v0/z2/z7/_036_ ;
 wire \v0/z2/z7/_037_ ;
 wire \v0/z2/z7/_038_ ;
 wire \v0/z2/z7/_039_ ;
 wire \v0/z2/z7/_040_ ;
 wire \v0/z2/z7/_041_ ;
 wire \v0/z2/z7/_042_ ;
 wire \v0/z2/z7/_043_ ;
 wire \v0/z2/z7/_044_ ;
 wire \v0/z2/z7/_045_ ;
 wire \v0/z2/z7/_046_ ;
 wire \v0/z2/z7/_047_ ;
 wire \v0/z2/z7/_048_ ;
 wire \v0/z2/z7/_049_ ;
 wire \v0/z3/_00_ ;
 wire \v0/z3/_01_ ;
 wire \v0/z3/_02_ ;
 wire \v0/z3/_03_ ;
 wire \v0/z3/_04_ ;
 wire \v0/z3/_05_ ;
 wire \v0/z3/_06_ ;
 wire \v0/z3/_07_ ;
 wire \v0/z3/_08_ ;
 wire \v0/z3/_09_ ;
 wire \v0/z3/_10_ ;
 wire \v0/z3/_11_ ;
 wire \v0/z3/_12_ ;
 wire \v0/z3/_13_ ;
 wire \v0/z3/_14_ ;
 wire \v0/z3/_15_ ;
 wire \v0/z3/_16_ ;
 wire \v0/z3/_17_ ;
 wire \v0/z3/_18_ ;
 wire \v0/z3/z1/_00_ ;
 wire \v0/z3/z1/_01_ ;
 wire \v0/z3/z1/_02_ ;
 wire \v0/z3/z1/_03_ ;
 wire \v0/z3/z1/_04_ ;
 wire \v0/z3/z1/_05_ ;
 wire \v0/z3/z1/_06_ ;
 wire \v0/z3/z1/_07_ ;
 wire \v0/z3/z1/_08_ ;
 wire \v0/z3/z1/_09_ ;
 wire \v0/z3/z1/_10_ ;
 wire \v0/z3/z1/z5/Cout ;
 wire \v0/z3/z1/z5/_00_ ;
 wire \v0/z3/z1/z5/_01_ ;
 wire \v0/z3/z1/z5/_02_ ;
 wire \v0/z3/z1/z5/_03_ ;
 wire \v0/z3/z1/z5/_04_ ;
 wire \v0/z3/z1/z5/_05_ ;
 wire \v0/z3/z1/z5/_06_ ;
 wire \v0/z3/z1/z6/Cout ;
 wire \v0/z3/z1/z6/_00_ ;
 wire \v0/z3/z1/z6/_01_ ;
 wire \v0/z3/z1/z6/_02_ ;
 wire \v0/z3/z1/z6/_03_ ;
 wire \v0/z3/z1/z6/_04_ ;
 wire \v0/z3/z1/z6/_05_ ;
 wire \v0/z3/z1/z6/_06_ ;
 wire \v0/z3/z1/z6/_07_ ;
 wire \v0/z3/z1/z6/_08_ ;
 wire \v0/z3/z1/z6/_09_ ;
 wire \v0/z3/z1/z6/_10_ ;
 wire \v0/z3/z1/z6/_11_ ;
 wire \v0/z3/z1/z6/_12_ ;
 wire \v0/z3/z1/z6/_13_ ;
 wire \v0/z3/z1/z6/_14_ ;
 wire \v0/z3/z1/z6/_15_ ;
 wire \v0/z3/z1/z6/_16_ ;
 wire \v0/z3/z1/z6/_17_ ;
 wire \v0/z3/z1/z6/_18_ ;
 wire \v0/z3/z1/z7/Cout ;
 wire \v0/z3/z1/z7/_00_ ;
 wire \v0/z3/z1/z7/_01_ ;
 wire \v0/z3/z1/z7/_02_ ;
 wire \v0/z3/z1/z7/_03_ ;
 wire \v0/z3/z1/z7/_04_ ;
 wire \v0/z3/z1/z7/_05_ ;
 wire \v0/z3/z1/z7/_06_ ;
 wire \v0/z3/z1/z7/_07_ ;
 wire \v0/z3/z1/z7/_08_ ;
 wire \v0/z3/z1/z7/_09_ ;
 wire \v0/z3/z1/z7/_10_ ;
 wire \v0/z3/z1/z7/_11_ ;
 wire \v0/z3/z1/z7/_12_ ;
 wire \v0/z3/z1/z7/_13_ ;
 wire \v0/z3/z1/z7/_14_ ;
 wire \v0/z3/z1/z7/_15_ ;
 wire \v0/z3/z1/z7/_16_ ;
 wire \v0/z3/z1/z7/_17_ ;
 wire \v0/z3/z1/z7/_18_ ;
 wire \v0/z3/z2/_00_ ;
 wire \v0/z3/z2/_01_ ;
 wire \v0/z3/z2/_02_ ;
 wire \v0/z3/z2/_03_ ;
 wire \v0/z3/z2/_04_ ;
 wire \v0/z3/z2/_05_ ;
 wire \v0/z3/z2/_06_ ;
 wire \v0/z3/z2/_07_ ;
 wire \v0/z3/z2/_08_ ;
 wire \v0/z3/z2/_09_ ;
 wire \v0/z3/z2/_10_ ;
 wire \v0/z3/z2/z5/Cout ;
 wire \v0/z3/z2/z5/_00_ ;
 wire \v0/z3/z2/z5/_01_ ;
 wire \v0/z3/z2/z5/_02_ ;
 wire \v0/z3/z2/z5/_03_ ;
 wire \v0/z3/z2/z5/_04_ ;
 wire \v0/z3/z2/z5/_05_ ;
 wire \v0/z3/z2/z5/_06_ ;
 wire \v0/z3/z2/z6/Cout ;
 wire \v0/z3/z2/z6/_00_ ;
 wire \v0/z3/z2/z6/_01_ ;
 wire \v0/z3/z2/z6/_02_ ;
 wire \v0/z3/z2/z6/_03_ ;
 wire \v0/z3/z2/z6/_04_ ;
 wire \v0/z3/z2/z6/_05_ ;
 wire \v0/z3/z2/z6/_06_ ;
 wire \v0/z3/z2/z6/_07_ ;
 wire \v0/z3/z2/z6/_08_ ;
 wire \v0/z3/z2/z6/_09_ ;
 wire \v0/z3/z2/z6/_10_ ;
 wire \v0/z3/z2/z6/_11_ ;
 wire \v0/z3/z2/z6/_12_ ;
 wire \v0/z3/z2/z6/_13_ ;
 wire \v0/z3/z2/z6/_14_ ;
 wire \v0/z3/z2/z6/_15_ ;
 wire \v0/z3/z2/z6/_16_ ;
 wire \v0/z3/z2/z6/_17_ ;
 wire \v0/z3/z2/z6/_18_ ;
 wire \v0/z3/z2/z7/Cout ;
 wire \v0/z3/z2/z7/_00_ ;
 wire \v0/z3/z2/z7/_01_ ;
 wire \v0/z3/z2/z7/_02_ ;
 wire \v0/z3/z2/z7/_03_ ;
 wire \v0/z3/z2/z7/_04_ ;
 wire \v0/z3/z2/z7/_05_ ;
 wire \v0/z3/z2/z7/_06_ ;
 wire \v0/z3/z2/z7/_07_ ;
 wire \v0/z3/z2/z7/_08_ ;
 wire \v0/z3/z2/z7/_09_ ;
 wire \v0/z3/z2/z7/_10_ ;
 wire \v0/z3/z2/z7/_11_ ;
 wire \v0/z3/z2/z7/_12_ ;
 wire \v0/z3/z2/z7/_13_ ;
 wire \v0/z3/z2/z7/_14_ ;
 wire \v0/z3/z2/z7/_15_ ;
 wire \v0/z3/z2/z7/_16_ ;
 wire \v0/z3/z2/z7/_17_ ;
 wire \v0/z3/z2/z7/_18_ ;
 wire \v0/z3/z3/_00_ ;
 wire \v0/z3/z3/_01_ ;
 wire \v0/z3/z3/_02_ ;
 wire \v0/z3/z3/_03_ ;
 wire \v0/z3/z3/_04_ ;
 wire \v0/z3/z3/_05_ ;
 wire \v0/z3/z3/_06_ ;
 wire \v0/z3/z3/_07_ ;
 wire \v0/z3/z3/_08_ ;
 wire \v0/z3/z3/_09_ ;
 wire \v0/z3/z3/_10_ ;
 wire \v0/z3/z3/z5/Cout ;
 wire \v0/z3/z3/z5/_00_ ;
 wire \v0/z3/z3/z5/_01_ ;
 wire \v0/z3/z3/z5/_02_ ;
 wire \v0/z3/z3/z5/_03_ ;
 wire \v0/z3/z3/z5/_04_ ;
 wire \v0/z3/z3/z5/_05_ ;
 wire \v0/z3/z3/z5/_06_ ;
 wire \v0/z3/z3/z6/Cout ;
 wire \v0/z3/z3/z6/_00_ ;
 wire \v0/z3/z3/z6/_01_ ;
 wire \v0/z3/z3/z6/_02_ ;
 wire \v0/z3/z3/z6/_03_ ;
 wire \v0/z3/z3/z6/_04_ ;
 wire \v0/z3/z3/z6/_05_ ;
 wire \v0/z3/z3/z6/_06_ ;
 wire \v0/z3/z3/z6/_07_ ;
 wire \v0/z3/z3/z6/_08_ ;
 wire \v0/z3/z3/z6/_09_ ;
 wire \v0/z3/z3/z6/_10_ ;
 wire \v0/z3/z3/z6/_11_ ;
 wire \v0/z3/z3/z6/_12_ ;
 wire \v0/z3/z3/z6/_13_ ;
 wire \v0/z3/z3/z6/_14_ ;
 wire \v0/z3/z3/z6/_15_ ;
 wire \v0/z3/z3/z6/_16_ ;
 wire \v0/z3/z3/z6/_17_ ;
 wire \v0/z3/z3/z6/_18_ ;
 wire \v0/z3/z3/z7/Cout ;
 wire \v0/z3/z3/z7/_00_ ;
 wire \v0/z3/z3/z7/_01_ ;
 wire \v0/z3/z3/z7/_02_ ;
 wire \v0/z3/z3/z7/_03_ ;
 wire \v0/z3/z3/z7/_04_ ;
 wire \v0/z3/z3/z7/_05_ ;
 wire \v0/z3/z3/z7/_06_ ;
 wire \v0/z3/z3/z7/_07_ ;
 wire \v0/z3/z3/z7/_08_ ;
 wire \v0/z3/z3/z7/_09_ ;
 wire \v0/z3/z3/z7/_10_ ;
 wire \v0/z3/z3/z7/_11_ ;
 wire \v0/z3/z3/z7/_12_ ;
 wire \v0/z3/z3/z7/_13_ ;
 wire \v0/z3/z3/z7/_14_ ;
 wire \v0/z3/z3/z7/_15_ ;
 wire \v0/z3/z3/z7/_16_ ;
 wire \v0/z3/z3/z7/_17_ ;
 wire \v0/z3/z3/z7/_18_ ;
 wire \v0/z3/z4/_00_ ;
 wire \v0/z3/z4/_01_ ;
 wire \v0/z3/z4/_02_ ;
 wire \v0/z3/z4/_03_ ;
 wire \v0/z3/z4/_04_ ;
 wire \v0/z3/z4/_05_ ;
 wire \v0/z3/z4/_06_ ;
 wire \v0/z3/z4/_07_ ;
 wire \v0/z3/z4/_08_ ;
 wire \v0/z3/z4/_09_ ;
 wire \v0/z3/z4/_10_ ;
 wire \v0/z3/z4/z5/Cout ;
 wire \v0/z3/z4/z5/_00_ ;
 wire \v0/z3/z4/z5/_01_ ;
 wire \v0/z3/z4/z5/_02_ ;
 wire \v0/z3/z4/z5/_03_ ;
 wire \v0/z3/z4/z5/_04_ ;
 wire \v0/z3/z4/z5/_05_ ;
 wire \v0/z3/z4/z5/_06_ ;
 wire \v0/z3/z4/z6/Cout ;
 wire \v0/z3/z4/z6/_00_ ;
 wire \v0/z3/z4/z6/_01_ ;
 wire \v0/z3/z4/z6/_02_ ;
 wire \v0/z3/z4/z6/_03_ ;
 wire \v0/z3/z4/z6/_04_ ;
 wire \v0/z3/z4/z6/_05_ ;
 wire \v0/z3/z4/z6/_06_ ;
 wire \v0/z3/z4/z6/_07_ ;
 wire \v0/z3/z4/z6/_08_ ;
 wire \v0/z3/z4/z6/_09_ ;
 wire \v0/z3/z4/z6/_10_ ;
 wire \v0/z3/z4/z6/_11_ ;
 wire \v0/z3/z4/z6/_12_ ;
 wire \v0/z3/z4/z6/_13_ ;
 wire \v0/z3/z4/z6/_14_ ;
 wire \v0/z3/z4/z6/_15_ ;
 wire \v0/z3/z4/z6/_16_ ;
 wire \v0/z3/z4/z6/_17_ ;
 wire \v0/z3/z4/z6/_18_ ;
 wire \v0/z3/z4/z7/Cout ;
 wire \v0/z3/z4/z7/_00_ ;
 wire \v0/z3/z4/z7/_01_ ;
 wire \v0/z3/z4/z7/_02_ ;
 wire \v0/z3/z4/z7/_03_ ;
 wire \v0/z3/z4/z7/_04_ ;
 wire \v0/z3/z4/z7/_05_ ;
 wire \v0/z3/z4/z7/_06_ ;
 wire \v0/z3/z4/z7/_07_ ;
 wire \v0/z3/z4/z7/_08_ ;
 wire \v0/z3/z4/z7/_09_ ;
 wire \v0/z3/z4/z7/_10_ ;
 wire \v0/z3/z4/z7/_11_ ;
 wire \v0/z3/z4/z7/_12_ ;
 wire \v0/z3/z4/z7/_13_ ;
 wire \v0/z3/z4/z7/_14_ ;
 wire \v0/z3/z4/z7/_15_ ;
 wire \v0/z3/z4/z7/_16_ ;
 wire \v0/z3/z4/z7/_17_ ;
 wire \v0/z3/z4/z7/_18_ ;
 wire \v0/z3/z5/Cout ;
 wire \v0/z3/z5/_00_ ;
 wire \v0/z3/z5/_01_ ;
 wire \v0/z3/z5/_02_ ;
 wire \v0/z3/z5/_03_ ;
 wire \v0/z3/z5/_04_ ;
 wire \v0/z3/z5/_05_ ;
 wire \v0/z3/z5/_06_ ;
 wire \v0/z3/z5/_07_ ;
 wire \v0/z3/z5/_08_ ;
 wire \v0/z3/z5/_09_ ;
 wire \v0/z3/z5/_10_ ;
 wire \v0/z3/z5/_11_ ;
 wire \v0/z3/z5/_12_ ;
 wire \v0/z3/z5/_13_ ;
 wire \v0/z3/z5/_14_ ;
 wire \v0/z3/z5/_15_ ;
 wire \v0/z3/z5/_16_ ;
 wire \v0/z3/z5/_17_ ;
 wire \v0/z3/z5/_18_ ;
 wire \v0/z3/z5/_19_ ;
 wire \v0/z3/z5/_20_ ;
 wire \v0/z3/z5/_21_ ;
 wire \v0/z3/z5/_22_ ;
 wire \v0/z3/z5/_23_ ;
 wire \v0/z3/z5/_24_ ;
 wire \v0/z3/z5/_25_ ;
 wire \v0/z3/z5/_26_ ;
 wire \v0/z3/z6/Cout ;
 wire \v0/z3/z6/_000_ ;
 wire \v0/z3/z6/_001_ ;
 wire \v0/z3/z6/_002_ ;
 wire \v0/z3/z6/_003_ ;
 wire \v0/z3/z6/_004_ ;
 wire \v0/z3/z6/_005_ ;
 wire \v0/z3/z6/_006_ ;
 wire \v0/z3/z6/_007_ ;
 wire \v0/z3/z6/_008_ ;
 wire \v0/z3/z6/_009_ ;
 wire \v0/z3/z6/_010_ ;
 wire \v0/z3/z6/_011_ ;
 wire \v0/z3/z6/_012_ ;
 wire \v0/z3/z6/_013_ ;
 wire \v0/z3/z6/_014_ ;
 wire \v0/z3/z6/_015_ ;
 wire \v0/z3/z6/_016_ ;
 wire \v0/z3/z6/_017_ ;
 wire \v0/z3/z6/_018_ ;
 wire \v0/z3/z6/_019_ ;
 wire \v0/z3/z6/_020_ ;
 wire \v0/z3/z6/_021_ ;
 wire \v0/z3/z6/_022_ ;
 wire \v0/z3/z6/_023_ ;
 wire \v0/z3/z6/_024_ ;
 wire \v0/z3/z6/_025_ ;
 wire \v0/z3/z6/_026_ ;
 wire \v0/z3/z6/_027_ ;
 wire \v0/z3/z6/_028_ ;
 wire \v0/z3/z6/_029_ ;
 wire \v0/z3/z6/_030_ ;
 wire \v0/z3/z6/_031_ ;
 wire \v0/z3/z6/_032_ ;
 wire \v0/z3/z6/_033_ ;
 wire \v0/z3/z6/_034_ ;
 wire \v0/z3/z6/_035_ ;
 wire \v0/z3/z6/_036_ ;
 wire \v0/z3/z6/_037_ ;
 wire \v0/z3/z6/_038_ ;
 wire \v0/z3/z6/_039_ ;
 wire \v0/z3/z6/_040_ ;
 wire \v0/z3/z6/_041_ ;
 wire \v0/z3/z6/_042_ ;
 wire \v0/z3/z6/_043_ ;
 wire \v0/z3/z6/_044_ ;
 wire \v0/z3/z6/_045_ ;
 wire \v0/z3/z6/_046_ ;
 wire \v0/z3/z6/_047_ ;
 wire \v0/z3/z6/_048_ ;
 wire \v0/z3/z6/_049_ ;
 wire \v0/z3/z7/Cout ;
 wire \v0/z3/z7/_000_ ;
 wire \v0/z3/z7/_001_ ;
 wire \v0/z3/z7/_002_ ;
 wire \v0/z3/z7/_003_ ;
 wire \v0/z3/z7/_004_ ;
 wire \v0/z3/z7/_005_ ;
 wire \v0/z3/z7/_006_ ;
 wire \v0/z3/z7/_007_ ;
 wire \v0/z3/z7/_008_ ;
 wire \v0/z3/z7/_009_ ;
 wire \v0/z3/z7/_010_ ;
 wire \v0/z3/z7/_011_ ;
 wire \v0/z3/z7/_012_ ;
 wire \v0/z3/z7/_013_ ;
 wire \v0/z3/z7/_014_ ;
 wire \v0/z3/z7/_015_ ;
 wire \v0/z3/z7/_016_ ;
 wire \v0/z3/z7/_017_ ;
 wire \v0/z3/z7/_018_ ;
 wire \v0/z3/z7/_019_ ;
 wire \v0/z3/z7/_020_ ;
 wire \v0/z3/z7/_021_ ;
 wire \v0/z3/z7/_022_ ;
 wire \v0/z3/z7/_023_ ;
 wire \v0/z3/z7/_024_ ;
 wire \v0/z3/z7/_025_ ;
 wire \v0/z3/z7/_026_ ;
 wire \v0/z3/z7/_027_ ;
 wire \v0/z3/z7/_028_ ;
 wire \v0/z3/z7/_029_ ;
 wire \v0/z3/z7/_030_ ;
 wire \v0/z3/z7/_031_ ;
 wire \v0/z3/z7/_032_ ;
 wire \v0/z3/z7/_033_ ;
 wire \v0/z3/z7/_034_ ;
 wire \v0/z3/z7/_035_ ;
 wire \v0/z3/z7/_036_ ;
 wire \v0/z3/z7/_037_ ;
 wire \v0/z3/z7/_038_ ;
 wire \v0/z3/z7/_039_ ;
 wire \v0/z3/z7/_040_ ;
 wire \v0/z3/z7/_041_ ;
 wire \v0/z3/z7/_042_ ;
 wire \v0/z3/z7/_043_ ;
 wire \v0/z3/z7/_044_ ;
 wire \v0/z3/z7/_045_ ;
 wire \v0/z3/z7/_046_ ;
 wire \v0/z3/z7/_047_ ;
 wire \v0/z3/z7/_048_ ;
 wire \v0/z3/z7/_049_ ;
 wire \v0/z4/_00_ ;
 wire \v0/z4/_01_ ;
 wire \v0/z4/_02_ ;
 wire \v0/z4/_03_ ;
 wire \v0/z4/_04_ ;
 wire \v0/z4/_05_ ;
 wire \v0/z4/_06_ ;
 wire \v0/z4/_07_ ;
 wire \v0/z4/_08_ ;
 wire \v0/z4/_09_ ;
 wire \v0/z4/_10_ ;
 wire \v0/z4/_11_ ;
 wire \v0/z4/_12_ ;
 wire \v0/z4/_13_ ;
 wire \v0/z4/_14_ ;
 wire \v0/z4/_15_ ;
 wire \v0/z4/_16_ ;
 wire \v0/z4/_17_ ;
 wire \v0/z4/_18_ ;
 wire \v0/z4/z1/_00_ ;
 wire \v0/z4/z1/_01_ ;
 wire \v0/z4/z1/_02_ ;
 wire \v0/z4/z1/_03_ ;
 wire \v0/z4/z1/_04_ ;
 wire \v0/z4/z1/_05_ ;
 wire \v0/z4/z1/_06_ ;
 wire \v0/z4/z1/_07_ ;
 wire \v0/z4/z1/_08_ ;
 wire \v0/z4/z1/_09_ ;
 wire \v0/z4/z1/_10_ ;
 wire \v0/z4/z1/z5/Cout ;
 wire \v0/z4/z1/z5/_00_ ;
 wire \v0/z4/z1/z5/_01_ ;
 wire \v0/z4/z1/z5/_02_ ;
 wire \v0/z4/z1/z5/_03_ ;
 wire \v0/z4/z1/z5/_04_ ;
 wire \v0/z4/z1/z5/_05_ ;
 wire \v0/z4/z1/z5/_06_ ;
 wire \v0/z4/z1/z6/Cout ;
 wire \v0/z4/z1/z6/_00_ ;
 wire \v0/z4/z1/z6/_01_ ;
 wire \v0/z4/z1/z6/_02_ ;
 wire \v0/z4/z1/z6/_03_ ;
 wire \v0/z4/z1/z6/_04_ ;
 wire \v0/z4/z1/z6/_05_ ;
 wire \v0/z4/z1/z6/_06_ ;
 wire \v0/z4/z1/z6/_07_ ;
 wire \v0/z4/z1/z6/_08_ ;
 wire \v0/z4/z1/z6/_09_ ;
 wire \v0/z4/z1/z6/_10_ ;
 wire \v0/z4/z1/z6/_11_ ;
 wire \v0/z4/z1/z6/_12_ ;
 wire \v0/z4/z1/z6/_13_ ;
 wire \v0/z4/z1/z6/_14_ ;
 wire \v0/z4/z1/z6/_15_ ;
 wire \v0/z4/z1/z6/_16_ ;
 wire \v0/z4/z1/z6/_17_ ;
 wire \v0/z4/z1/z6/_18_ ;
 wire \v0/z4/z1/z7/Cout ;
 wire \v0/z4/z1/z7/_00_ ;
 wire \v0/z4/z1/z7/_01_ ;
 wire \v0/z4/z1/z7/_02_ ;
 wire \v0/z4/z1/z7/_03_ ;
 wire \v0/z4/z1/z7/_04_ ;
 wire \v0/z4/z1/z7/_05_ ;
 wire \v0/z4/z1/z7/_06_ ;
 wire \v0/z4/z1/z7/_07_ ;
 wire \v0/z4/z1/z7/_08_ ;
 wire \v0/z4/z1/z7/_09_ ;
 wire \v0/z4/z1/z7/_10_ ;
 wire \v0/z4/z1/z7/_11_ ;
 wire \v0/z4/z1/z7/_12_ ;
 wire \v0/z4/z1/z7/_13_ ;
 wire \v0/z4/z1/z7/_14_ ;
 wire \v0/z4/z1/z7/_15_ ;
 wire \v0/z4/z1/z7/_16_ ;
 wire \v0/z4/z1/z7/_17_ ;
 wire \v0/z4/z1/z7/_18_ ;
 wire \v0/z4/z2/_00_ ;
 wire \v0/z4/z2/_01_ ;
 wire \v0/z4/z2/_02_ ;
 wire \v0/z4/z2/_03_ ;
 wire \v0/z4/z2/_04_ ;
 wire \v0/z4/z2/_05_ ;
 wire \v0/z4/z2/_06_ ;
 wire \v0/z4/z2/_07_ ;
 wire \v0/z4/z2/_08_ ;
 wire \v0/z4/z2/_09_ ;
 wire \v0/z4/z2/_10_ ;
 wire \v0/z4/z2/z5/Cout ;
 wire \v0/z4/z2/z5/_00_ ;
 wire \v0/z4/z2/z5/_01_ ;
 wire \v0/z4/z2/z5/_02_ ;
 wire \v0/z4/z2/z5/_03_ ;
 wire \v0/z4/z2/z5/_04_ ;
 wire \v0/z4/z2/z5/_05_ ;
 wire \v0/z4/z2/z5/_06_ ;
 wire \v0/z4/z2/z6/Cout ;
 wire \v0/z4/z2/z6/_00_ ;
 wire \v0/z4/z2/z6/_01_ ;
 wire \v0/z4/z2/z6/_02_ ;
 wire \v0/z4/z2/z6/_03_ ;
 wire \v0/z4/z2/z6/_04_ ;
 wire \v0/z4/z2/z6/_05_ ;
 wire \v0/z4/z2/z6/_06_ ;
 wire \v0/z4/z2/z6/_07_ ;
 wire \v0/z4/z2/z6/_08_ ;
 wire \v0/z4/z2/z6/_09_ ;
 wire \v0/z4/z2/z6/_10_ ;
 wire \v0/z4/z2/z6/_11_ ;
 wire \v0/z4/z2/z6/_12_ ;
 wire \v0/z4/z2/z6/_13_ ;
 wire \v0/z4/z2/z6/_14_ ;
 wire \v0/z4/z2/z6/_15_ ;
 wire \v0/z4/z2/z6/_16_ ;
 wire \v0/z4/z2/z6/_17_ ;
 wire \v0/z4/z2/z6/_18_ ;
 wire \v0/z4/z2/z7/Cout ;
 wire \v0/z4/z2/z7/_00_ ;
 wire \v0/z4/z2/z7/_01_ ;
 wire \v0/z4/z2/z7/_02_ ;
 wire \v0/z4/z2/z7/_03_ ;
 wire \v0/z4/z2/z7/_04_ ;
 wire \v0/z4/z2/z7/_05_ ;
 wire \v0/z4/z2/z7/_06_ ;
 wire \v0/z4/z2/z7/_07_ ;
 wire \v0/z4/z2/z7/_08_ ;
 wire \v0/z4/z2/z7/_09_ ;
 wire \v0/z4/z2/z7/_10_ ;
 wire \v0/z4/z2/z7/_11_ ;
 wire \v0/z4/z2/z7/_12_ ;
 wire \v0/z4/z2/z7/_13_ ;
 wire \v0/z4/z2/z7/_14_ ;
 wire \v0/z4/z2/z7/_15_ ;
 wire \v0/z4/z2/z7/_16_ ;
 wire \v0/z4/z2/z7/_17_ ;
 wire \v0/z4/z2/z7/_18_ ;
 wire \v0/z4/z3/_00_ ;
 wire \v0/z4/z3/_01_ ;
 wire \v0/z4/z3/_02_ ;
 wire \v0/z4/z3/_03_ ;
 wire \v0/z4/z3/_04_ ;
 wire \v0/z4/z3/_05_ ;
 wire \v0/z4/z3/_06_ ;
 wire \v0/z4/z3/_07_ ;
 wire \v0/z4/z3/_08_ ;
 wire \v0/z4/z3/_09_ ;
 wire \v0/z4/z3/_10_ ;
 wire \v0/z4/z3/z5/Cout ;
 wire \v0/z4/z3/z5/_00_ ;
 wire \v0/z4/z3/z5/_01_ ;
 wire \v0/z4/z3/z5/_02_ ;
 wire \v0/z4/z3/z5/_03_ ;
 wire \v0/z4/z3/z5/_04_ ;
 wire \v0/z4/z3/z5/_05_ ;
 wire \v0/z4/z3/z5/_06_ ;
 wire \v0/z4/z3/z6/Cout ;
 wire \v0/z4/z3/z6/_00_ ;
 wire \v0/z4/z3/z6/_01_ ;
 wire \v0/z4/z3/z6/_02_ ;
 wire \v0/z4/z3/z6/_03_ ;
 wire \v0/z4/z3/z6/_04_ ;
 wire \v0/z4/z3/z6/_05_ ;
 wire \v0/z4/z3/z6/_06_ ;
 wire \v0/z4/z3/z6/_07_ ;
 wire \v0/z4/z3/z6/_08_ ;
 wire \v0/z4/z3/z6/_09_ ;
 wire \v0/z4/z3/z6/_10_ ;
 wire \v0/z4/z3/z6/_11_ ;
 wire \v0/z4/z3/z6/_12_ ;
 wire \v0/z4/z3/z6/_13_ ;
 wire \v0/z4/z3/z6/_14_ ;
 wire \v0/z4/z3/z6/_15_ ;
 wire \v0/z4/z3/z6/_16_ ;
 wire \v0/z4/z3/z6/_17_ ;
 wire \v0/z4/z3/z6/_18_ ;
 wire \v0/z4/z3/z7/Cout ;
 wire \v0/z4/z3/z7/_00_ ;
 wire \v0/z4/z3/z7/_01_ ;
 wire \v0/z4/z3/z7/_02_ ;
 wire \v0/z4/z3/z7/_03_ ;
 wire \v0/z4/z3/z7/_04_ ;
 wire \v0/z4/z3/z7/_05_ ;
 wire \v0/z4/z3/z7/_06_ ;
 wire \v0/z4/z3/z7/_07_ ;
 wire \v0/z4/z3/z7/_08_ ;
 wire \v0/z4/z3/z7/_09_ ;
 wire \v0/z4/z3/z7/_10_ ;
 wire \v0/z4/z3/z7/_11_ ;
 wire \v0/z4/z3/z7/_12_ ;
 wire \v0/z4/z3/z7/_13_ ;
 wire \v0/z4/z3/z7/_14_ ;
 wire \v0/z4/z3/z7/_15_ ;
 wire \v0/z4/z3/z7/_16_ ;
 wire \v0/z4/z3/z7/_17_ ;
 wire \v0/z4/z3/z7/_18_ ;
 wire \v0/z4/z4/_00_ ;
 wire \v0/z4/z4/_01_ ;
 wire \v0/z4/z4/_02_ ;
 wire \v0/z4/z4/_03_ ;
 wire \v0/z4/z4/_04_ ;
 wire \v0/z4/z4/_05_ ;
 wire \v0/z4/z4/_06_ ;
 wire \v0/z4/z4/_07_ ;
 wire \v0/z4/z4/_08_ ;
 wire \v0/z4/z4/_09_ ;
 wire \v0/z4/z4/_10_ ;
 wire \v0/z4/z4/z5/Cout ;
 wire \v0/z4/z4/z5/_00_ ;
 wire \v0/z4/z4/z5/_01_ ;
 wire \v0/z4/z4/z5/_02_ ;
 wire \v0/z4/z4/z5/_03_ ;
 wire \v0/z4/z4/z5/_04_ ;
 wire \v0/z4/z4/z5/_05_ ;
 wire \v0/z4/z4/z5/_06_ ;
 wire \v0/z4/z4/z6/Cout ;
 wire \v0/z4/z4/z6/_00_ ;
 wire \v0/z4/z4/z6/_01_ ;
 wire \v0/z4/z4/z6/_02_ ;
 wire \v0/z4/z4/z6/_03_ ;
 wire \v0/z4/z4/z6/_04_ ;
 wire \v0/z4/z4/z6/_05_ ;
 wire \v0/z4/z4/z6/_06_ ;
 wire \v0/z4/z4/z6/_07_ ;
 wire \v0/z4/z4/z6/_08_ ;
 wire \v0/z4/z4/z6/_09_ ;
 wire \v0/z4/z4/z6/_10_ ;
 wire \v0/z4/z4/z6/_11_ ;
 wire \v0/z4/z4/z6/_12_ ;
 wire \v0/z4/z4/z6/_13_ ;
 wire \v0/z4/z4/z6/_14_ ;
 wire \v0/z4/z4/z6/_15_ ;
 wire \v0/z4/z4/z6/_16_ ;
 wire \v0/z4/z4/z6/_17_ ;
 wire \v0/z4/z4/z6/_18_ ;
 wire \v0/z4/z4/z7/Cout ;
 wire \v0/z4/z4/z7/_00_ ;
 wire \v0/z4/z4/z7/_01_ ;
 wire \v0/z4/z4/z7/_02_ ;
 wire \v0/z4/z4/z7/_03_ ;
 wire \v0/z4/z4/z7/_04_ ;
 wire \v0/z4/z4/z7/_05_ ;
 wire \v0/z4/z4/z7/_06_ ;
 wire \v0/z4/z4/z7/_07_ ;
 wire \v0/z4/z4/z7/_08_ ;
 wire \v0/z4/z4/z7/_09_ ;
 wire \v0/z4/z4/z7/_10_ ;
 wire \v0/z4/z4/z7/_11_ ;
 wire \v0/z4/z4/z7/_12_ ;
 wire \v0/z4/z4/z7/_13_ ;
 wire \v0/z4/z4/z7/_14_ ;
 wire \v0/z4/z4/z7/_15_ ;
 wire \v0/z4/z4/z7/_16_ ;
 wire \v0/z4/z4/z7/_17_ ;
 wire \v0/z4/z4/z7/_18_ ;
 wire \v0/z4/z5/Cout ;
 wire \v0/z4/z5/_00_ ;
 wire \v0/z4/z5/_01_ ;
 wire \v0/z4/z5/_02_ ;
 wire \v0/z4/z5/_03_ ;
 wire \v0/z4/z5/_04_ ;
 wire \v0/z4/z5/_05_ ;
 wire \v0/z4/z5/_06_ ;
 wire \v0/z4/z5/_07_ ;
 wire \v0/z4/z5/_08_ ;
 wire \v0/z4/z5/_09_ ;
 wire \v0/z4/z5/_10_ ;
 wire \v0/z4/z5/_11_ ;
 wire \v0/z4/z5/_12_ ;
 wire \v0/z4/z5/_13_ ;
 wire \v0/z4/z5/_14_ ;
 wire \v0/z4/z5/_15_ ;
 wire \v0/z4/z5/_16_ ;
 wire \v0/z4/z5/_17_ ;
 wire \v0/z4/z5/_18_ ;
 wire \v0/z4/z5/_19_ ;
 wire \v0/z4/z5/_20_ ;
 wire \v0/z4/z5/_21_ ;
 wire \v0/z4/z5/_22_ ;
 wire \v0/z4/z5/_23_ ;
 wire \v0/z4/z5/_24_ ;
 wire \v0/z4/z5/_25_ ;
 wire \v0/z4/z5/_26_ ;
 wire \v0/z4/z6/Cout ;
 wire \v0/z4/z6/_000_ ;
 wire \v0/z4/z6/_001_ ;
 wire \v0/z4/z6/_002_ ;
 wire \v0/z4/z6/_003_ ;
 wire \v0/z4/z6/_004_ ;
 wire \v0/z4/z6/_005_ ;
 wire \v0/z4/z6/_006_ ;
 wire \v0/z4/z6/_007_ ;
 wire \v0/z4/z6/_008_ ;
 wire \v0/z4/z6/_009_ ;
 wire \v0/z4/z6/_010_ ;
 wire \v0/z4/z6/_011_ ;
 wire \v0/z4/z6/_012_ ;
 wire \v0/z4/z6/_013_ ;
 wire \v0/z4/z6/_014_ ;
 wire \v0/z4/z6/_015_ ;
 wire \v0/z4/z6/_016_ ;
 wire \v0/z4/z6/_017_ ;
 wire \v0/z4/z6/_018_ ;
 wire \v0/z4/z6/_019_ ;
 wire \v0/z4/z6/_020_ ;
 wire \v0/z4/z6/_021_ ;
 wire \v0/z4/z6/_022_ ;
 wire \v0/z4/z6/_023_ ;
 wire \v0/z4/z6/_024_ ;
 wire \v0/z4/z6/_025_ ;
 wire \v0/z4/z6/_026_ ;
 wire \v0/z4/z6/_027_ ;
 wire \v0/z4/z6/_028_ ;
 wire \v0/z4/z6/_029_ ;
 wire \v0/z4/z6/_030_ ;
 wire \v0/z4/z6/_031_ ;
 wire \v0/z4/z6/_032_ ;
 wire \v0/z4/z6/_033_ ;
 wire \v0/z4/z6/_034_ ;
 wire \v0/z4/z6/_035_ ;
 wire \v0/z4/z6/_036_ ;
 wire \v0/z4/z6/_037_ ;
 wire \v0/z4/z6/_038_ ;
 wire \v0/z4/z6/_039_ ;
 wire \v0/z4/z6/_040_ ;
 wire \v0/z4/z6/_041_ ;
 wire \v0/z4/z6/_042_ ;
 wire \v0/z4/z6/_043_ ;
 wire \v0/z4/z6/_044_ ;
 wire \v0/z4/z6/_045_ ;
 wire \v0/z4/z6/_046_ ;
 wire \v0/z4/z6/_047_ ;
 wire \v0/z4/z6/_048_ ;
 wire \v0/z4/z6/_049_ ;
 wire \v0/z4/z7/Cout ;
 wire \v0/z4/z7/_000_ ;
 wire \v0/z4/z7/_001_ ;
 wire \v0/z4/z7/_002_ ;
 wire \v0/z4/z7/_003_ ;
 wire \v0/z4/z7/_004_ ;
 wire \v0/z4/z7/_005_ ;
 wire \v0/z4/z7/_006_ ;
 wire \v0/z4/z7/_007_ ;
 wire \v0/z4/z7/_008_ ;
 wire \v0/z4/z7/_009_ ;
 wire \v0/z4/z7/_010_ ;
 wire \v0/z4/z7/_011_ ;
 wire \v0/z4/z7/_012_ ;
 wire \v0/z4/z7/_013_ ;
 wire \v0/z4/z7/_014_ ;
 wire \v0/z4/z7/_015_ ;
 wire \v0/z4/z7/_016_ ;
 wire \v0/z4/z7/_017_ ;
 wire \v0/z4/z7/_018_ ;
 wire \v0/z4/z7/_019_ ;
 wire \v0/z4/z7/_020_ ;
 wire \v0/z4/z7/_021_ ;
 wire \v0/z4/z7/_022_ ;
 wire \v0/z4/z7/_023_ ;
 wire \v0/z4/z7/_024_ ;
 wire \v0/z4/z7/_025_ ;
 wire \v0/z4/z7/_026_ ;
 wire \v0/z4/z7/_027_ ;
 wire \v0/z4/z7/_028_ ;
 wire \v0/z4/z7/_029_ ;
 wire \v0/z4/z7/_030_ ;
 wire \v0/z4/z7/_031_ ;
 wire \v0/z4/z7/_032_ ;
 wire \v0/z4/z7/_033_ ;
 wire \v0/z4/z7/_034_ ;
 wire \v0/z4/z7/_035_ ;
 wire \v0/z4/z7/_036_ ;
 wire \v0/z4/z7/_037_ ;
 wire \v0/z4/z7/_038_ ;
 wire \v0/z4/z7/_039_ ;
 wire \v0/z4/z7/_040_ ;
 wire \v0/z4/z7/_041_ ;
 wire \v0/z4/z7/_042_ ;
 wire \v0/z4/z7/_043_ ;
 wire \v0/z4/z7/_044_ ;
 wire \v0/z4/z7/_045_ ;
 wire \v0/z4/z7/_046_ ;
 wire \v0/z4/z7/_047_ ;
 wire \v0/z4/z7/_048_ ;
 wire \v0/z4/z7/_049_ ;
 wire \v0/z5/Cout ;
 wire \v0/z5/_000_ ;
 wire \v0/z5/_001_ ;
 wire \v0/z5/_002_ ;
 wire \v0/z5/_003_ ;
 wire \v0/z5/_004_ ;
 wire \v0/z5/_005_ ;
 wire \v0/z5/_006_ ;
 wire \v0/z5/_007_ ;
 wire \v0/z5/_008_ ;
 wire \v0/z5/_009_ ;
 wire \v0/z5/_010_ ;
 wire \v0/z5/_011_ ;
 wire \v0/z5/_012_ ;
 wire \v0/z5/_013_ ;
 wire \v0/z5/_014_ ;
 wire \v0/z5/_015_ ;
 wire \v0/z5/_016_ ;
 wire \v0/z5/_017_ ;
 wire \v0/z5/_018_ ;
 wire \v0/z5/_019_ ;
 wire \v0/z5/_020_ ;
 wire \v0/z5/_021_ ;
 wire \v0/z5/_022_ ;
 wire \v0/z5/_023_ ;
 wire \v0/z5/_024_ ;
 wire \v0/z5/_025_ ;
 wire \v0/z5/_026_ ;
 wire \v0/z5/_027_ ;
 wire \v0/z5/_028_ ;
 wire \v0/z5/_029_ ;
 wire \v0/z5/_030_ ;
 wire \v0/z5/_031_ ;
 wire \v0/z5/_032_ ;
 wire \v0/z5/_033_ ;
 wire \v0/z5/_034_ ;
 wire \v0/z5/_035_ ;
 wire \v0/z5/_036_ ;
 wire \v0/z5/_037_ ;
 wire \v0/z5/_038_ ;
 wire \v0/z5/_039_ ;
 wire \v0/z5/_040_ ;
 wire \v0/z5/_041_ ;
 wire \v0/z5/_042_ ;
 wire \v0/z5/_043_ ;
 wire \v0/z5/_044_ ;
 wire \v0/z5/_045_ ;
 wire \v0/z5/_046_ ;
 wire \v0/z5/_047_ ;
 wire \v0/z5/_048_ ;
 wire \v0/z5/_049_ ;
 wire \v0/z5/_050_ ;
 wire \v0/z5/_051_ ;
 wire \v0/z5/_052_ ;
 wire \v0/z5/_053_ ;
 wire \v0/z5/_054_ ;
 wire \v0/z5/_055_ ;
 wire \v0/z5/_056_ ;
 wire \v0/z5/_057_ ;
 wire \v0/z5/_058_ ;
 wire \v0/z5/_059_ ;
 wire \v0/z5/_060_ ;
 wire \v0/z5/_061_ ;
 wire \v0/z5/_062_ ;
 wire \v0/z5/_063_ ;
 wire \v0/z5/_064_ ;
 wire \v0/z5/_065_ ;
 wire \v0/z5/_066_ ;
 wire \v0/z5/_067_ ;
 wire \v0/z5/_068_ ;
 wire \v0/z5/_069_ ;
 wire \v0/z6/Cout ;
 wire \v0/z6/_000_ ;
 wire \v0/z6/_001_ ;
 wire \v0/z6/_002_ ;
 wire \v0/z6/_003_ ;
 wire \v0/z6/_004_ ;
 wire \v0/z6/_005_ ;
 wire \v0/z6/_006_ ;
 wire \v0/z6/_007_ ;
 wire \v0/z6/_008_ ;
 wire \v0/z6/_009_ ;
 wire \v0/z6/_010_ ;
 wire \v0/z6/_011_ ;
 wire \v0/z6/_012_ ;
 wire \v0/z6/_013_ ;
 wire \v0/z6/_014_ ;
 wire \v0/z6/_015_ ;
 wire \v0/z6/_016_ ;
 wire \v0/z6/_017_ ;
 wire \v0/z6/_018_ ;
 wire \v0/z6/_019_ ;
 wire \v0/z6/_020_ ;
 wire \v0/z6/_021_ ;
 wire \v0/z6/_022_ ;
 wire \v0/z6/_023_ ;
 wire \v0/z6/_024_ ;
 wire \v0/z6/_025_ ;
 wire \v0/z6/_026_ ;
 wire \v0/z6/_027_ ;
 wire \v0/z6/_028_ ;
 wire \v0/z6/_029_ ;
 wire \v0/z6/_030_ ;
 wire \v0/z6/_031_ ;
 wire \v0/z6/_032_ ;
 wire \v0/z6/_033_ ;
 wire \v0/z6/_034_ ;
 wire \v0/z6/_035_ ;
 wire \v0/z6/_036_ ;
 wire \v0/z6/_037_ ;
 wire \v0/z6/_038_ ;
 wire \v0/z6/_039_ ;
 wire \v0/z6/_040_ ;
 wire \v0/z6/_041_ ;
 wire \v0/z6/_042_ ;
 wire \v0/z6/_043_ ;
 wire \v0/z6/_044_ ;
 wire \v0/z6/_045_ ;
 wire \v0/z6/_046_ ;
 wire \v0/z6/_047_ ;
 wire \v0/z6/_048_ ;
 wire \v0/z6/_049_ ;
 wire \v0/z6/_050_ ;
 wire \v0/z6/_051_ ;
 wire \v0/z6/_052_ ;
 wire \v0/z6/_053_ ;
 wire \v0/z6/_054_ ;
 wire \v0/z6/_055_ ;
 wire \v0/z6/_056_ ;
 wire \v0/z6/_057_ ;
 wire \v0/z6/_058_ ;
 wire \v0/z6/_059_ ;
 wire \v0/z6/_060_ ;
 wire \v0/z6/_061_ ;
 wire \v0/z6/_062_ ;
 wire \v0/z6/_063_ ;
 wire \v0/z6/_064_ ;
 wire \v0/z6/_065_ ;
 wire \v0/z6/_066_ ;
 wire \v0/z6/_067_ ;
 wire \v0/z6/_068_ ;
 wire \v0/z6/_069_ ;
 wire \v0/z6/_070_ ;
 wire \v0/z6/_071_ ;
 wire \v0/z6/_072_ ;
 wire \v0/z6/_073_ ;
 wire \v0/z6/_074_ ;
 wire \v0/z6/_075_ ;
 wire \v0/z6/_076_ ;
 wire \v0/z6/_077_ ;
 wire \v0/z6/_078_ ;
 wire \v0/z6/_079_ ;
 wire \v0/z6/_080_ ;
 wire \v0/z6/_081_ ;
 wire \v0/z6/_082_ ;
 wire \v0/z6/_083_ ;
 wire \v0/z6/_084_ ;
 wire \v0/z6/_085_ ;
 wire \v0/z6/_086_ ;
 wire \v0/z6/_087_ ;
 wire \v0/z6/_088_ ;
 wire \v0/z6/_089_ ;
 wire \v0/z6/_090_ ;
 wire \v0/z6/_091_ ;
 wire \v0/z6/_092_ ;
 wire \v0/z6/_093_ ;
 wire \v0/z6/_094_ ;
 wire \v0/z6/_095_ ;
 wire \v0/z6/_096_ ;
 wire \v0/z6/_097_ ;
 wire \v0/z6/_098_ ;
 wire \v0/z6/_099_ ;
 wire \v0/z6/_100_ ;
 wire \v0/z6/_101_ ;
 wire \v0/z6/_102_ ;
 wire \v0/z6/_103_ ;
 wire \v0/z6/_104_ ;
 wire \v0/z6/_105_ ;
 wire \v0/z6/_106_ ;
 wire \v0/z6/_107_ ;
 wire \v0/z6/_108_ ;
 wire \v0/z6/_109_ ;
 wire \v0/z6/_110_ ;
 wire \v0/z6/_111_ ;
 wire \v0/z6/_112_ ;
 wire \v0/z7/Cout ;
 wire \v0/z7/_000_ ;
 wire \v0/z7/_001_ ;
 wire \v0/z7/_002_ ;
 wire \v0/z7/_003_ ;
 wire \v0/z7/_004_ ;
 wire \v0/z7/_005_ ;
 wire \v0/z7/_006_ ;
 wire \v0/z7/_007_ ;
 wire \v0/z7/_008_ ;
 wire \v0/z7/_009_ ;
 wire \v0/z7/_010_ ;
 wire \v0/z7/_011_ ;
 wire \v0/z7/_012_ ;
 wire \v0/z7/_013_ ;
 wire \v0/z7/_014_ ;
 wire \v0/z7/_015_ ;
 wire \v0/z7/_016_ ;
 wire \v0/z7/_017_ ;
 wire \v0/z7/_018_ ;
 wire \v0/z7/_019_ ;
 wire \v0/z7/_020_ ;
 wire \v0/z7/_021_ ;
 wire \v0/z7/_022_ ;
 wire \v0/z7/_023_ ;
 wire \v0/z7/_024_ ;
 wire \v0/z7/_025_ ;
 wire \v0/z7/_026_ ;
 wire \v0/z7/_027_ ;
 wire \v0/z7/_028_ ;
 wire \v0/z7/_029_ ;
 wire \v0/z7/_030_ ;
 wire \v0/z7/_031_ ;
 wire \v0/z7/_032_ ;
 wire \v0/z7/_033_ ;
 wire \v0/z7/_034_ ;
 wire \v0/z7/_035_ ;
 wire \v0/z7/_036_ ;
 wire \v0/z7/_037_ ;
 wire \v0/z7/_038_ ;
 wire \v0/z7/_039_ ;
 wire \v0/z7/_040_ ;
 wire \v0/z7/_041_ ;
 wire \v0/z7/_042_ ;
 wire \v0/z7/_043_ ;
 wire \v0/z7/_044_ ;
 wire \v0/z7/_045_ ;
 wire \v0/z7/_046_ ;
 wire \v0/z7/_047_ ;
 wire \v0/z7/_048_ ;
 wire \v0/z7/_049_ ;
 wire \v0/z7/_050_ ;
 wire \v0/z7/_051_ ;
 wire \v0/z7/_052_ ;
 wire \v0/z7/_053_ ;
 wire \v0/z7/_054_ ;
 wire \v0/z7/_055_ ;
 wire \v0/z7/_056_ ;
 wire \v0/z7/_057_ ;
 wire \v0/z7/_058_ ;
 wire \v0/z7/_059_ ;
 wire \v0/z7/_060_ ;
 wire \v0/z7/_061_ ;
 wire \v0/z7/_062_ ;
 wire \v0/z7/_063_ ;
 wire \v0/z7/_064_ ;
 wire \v0/z7/_065_ ;
 wire \v0/z7/_066_ ;
 wire \v0/z7/_067_ ;
 wire \v0/z7/_068_ ;
 wire \v0/z7/_069_ ;
 wire \v0/z7/_070_ ;
 wire \v0/z7/_071_ ;
 wire \v0/z7/_072_ ;
 wire \v0/z7/_073_ ;
 wire \v0/z7/_074_ ;
 wire \v0/z7/_075_ ;
 wire \v0/z7/_076_ ;
 wire \v0/z7/_077_ ;
 wire \v0/z7/_078_ ;
 wire \v0/z7/_079_ ;
 wire \v0/z7/_080_ ;
 wire \v0/z7/_081_ ;
 wire \v0/z7/_082_ ;
 wire \v0/z7/_083_ ;
 wire \v0/z7/_084_ ;
 wire \v0/z7/_085_ ;
 wire \v0/z7/_086_ ;
 wire \v0/z7/_087_ ;
 wire \v0/z7/_088_ ;
 wire \v0/z7/_089_ ;
 wire \v0/z7/_090_ ;
 wire \v0/z7/_091_ ;
 wire \v0/z7/_092_ ;
 wire \v0/z7/_093_ ;
 wire \v0/z7/_094_ ;
 wire \v0/z7/_095_ ;
 wire \v0/z7/_096_ ;
 wire \v0/z7/_097_ ;
 wire \v0/z7/_098_ ;
 wire \v0/z7/_099_ ;
 wire \v0/z7/_100_ ;
 wire \v0/z7/_101_ ;
 wire \v0/z7/_102_ ;
 wire \v0/z7/_103_ ;
 wire \v0/z7/_104_ ;
 wire \v0/z7/_105_ ;
 wire \v0/z7/_106_ ;
 wire \v0/z7/_107_ ;
 wire \v0/z7/_108_ ;
 wire \v0/z7/_109_ ;
 wire \v0/z7/_110_ ;
 wire \v0/z7/_111_ ;
 wire \v0/z7/_112_ ;
 wire [15:0] abs_a;
 wire [15:0] abs_b;
 wire [31:0] nextinp;
 wire [31:0] unsign;
 wire [15:0] \v0/q0 ;
 wire [15:0] \v0/q1 ;
 wire [15:0] \v0/q2 ;
 wire [15:0] \v0/q3 ;
 wire [15:0] \v0/q4 ;
 wire [23:0] \v0/q5 ;
 wire [7:0] \v0/z1/q0 ;
 wire [7:0] \v0/z1/q1 ;
 wire [7:0] \v0/z1/q2 ;
 wire [7:0] \v0/z1/q3 ;
 wire [7:0] \v0/z1/q4 ;
 wire [11:0] \v0/z1/q5 ;
 wire [3:0] \v0/z1/z1/q0 ;
 wire [3:0] \v0/z1/z1/q1 ;
 wire [3:0] \v0/z1/z1/q2 ;
 wire [3:0] \v0/z1/z1/q3 ;
 wire [3:0] \v0/z1/z1/q4 ;
 wire [5:0] \v0/z1/z1/q5 ;
 wire [3:0] \v0/z1/z1/z1/temp ;
 wire [3:0] \v0/z1/z1/z2/temp ;
 wire [3:0] \v0/z1/z1/z3/temp ;
 wire [3:0] \v0/z1/z1/z4/temp ;
 wire [3:0] \v0/z1/z2/q0 ;
 wire [3:0] \v0/z1/z2/q1 ;
 wire [3:0] \v0/z1/z2/q2 ;
 wire [3:0] \v0/z1/z2/q3 ;
 wire [3:0] \v0/z1/z2/q4 ;
 wire [5:0] \v0/z1/z2/q5 ;
 wire [3:0] \v0/z1/z2/z1/temp ;
 wire [3:0] \v0/z1/z2/z2/temp ;
 wire [3:0] \v0/z1/z2/z3/temp ;
 wire [3:0] \v0/z1/z2/z4/temp ;
 wire [3:0] \v0/z1/z3/q0 ;
 wire [3:0] \v0/z1/z3/q1 ;
 wire [3:0] \v0/z1/z3/q2 ;
 wire [3:0] \v0/z1/z3/q3 ;
 wire [3:0] \v0/z1/z3/q4 ;
 wire [5:0] \v0/z1/z3/q5 ;
 wire [3:0] \v0/z1/z3/z1/temp ;
 wire [3:0] \v0/z1/z3/z2/temp ;
 wire [3:0] \v0/z1/z3/z3/temp ;
 wire [3:0] \v0/z1/z3/z4/temp ;
 wire [3:0] \v0/z1/z4/q0 ;
 wire [3:0] \v0/z1/z4/q1 ;
 wire [3:0] \v0/z1/z4/q2 ;
 wire [3:0] \v0/z1/z4/q3 ;
 wire [3:0] \v0/z1/z4/q4 ;
 wire [5:0] \v0/z1/z4/q5 ;
 wire [3:0] \v0/z1/z4/z1/temp ;
 wire [3:0] \v0/z1/z4/z2/temp ;
 wire [3:0] \v0/z1/z4/z3/temp ;
 wire [3:0] \v0/z1/z4/z4/temp ;
 wire [7:0] \v0/z2/q0 ;
 wire [7:0] \v0/z2/q1 ;
 wire [7:0] \v0/z2/q2 ;
 wire [7:0] \v0/z2/q3 ;
 wire [7:0] \v0/z2/q4 ;
 wire [11:0] \v0/z2/q5 ;
 wire [3:0] \v0/z2/z1/q0 ;
 wire [3:0] \v0/z2/z1/q1 ;
 wire [3:0] \v0/z2/z1/q2 ;
 wire [3:0] \v0/z2/z1/q3 ;
 wire [3:0] \v0/z2/z1/q4 ;
 wire [5:0] \v0/z2/z1/q5 ;
 wire [3:0] \v0/z2/z1/z1/temp ;
 wire [3:0] \v0/z2/z1/z2/temp ;
 wire [3:0] \v0/z2/z1/z3/temp ;
 wire [3:0] \v0/z2/z1/z4/temp ;
 wire [3:0] \v0/z2/z2/q0 ;
 wire [3:0] \v0/z2/z2/q1 ;
 wire [3:0] \v0/z2/z2/q2 ;
 wire [3:0] \v0/z2/z2/q3 ;
 wire [3:0] \v0/z2/z2/q4 ;
 wire [5:0] \v0/z2/z2/q5 ;
 wire [3:0] \v0/z2/z2/z1/temp ;
 wire [3:0] \v0/z2/z2/z2/temp ;
 wire [3:0] \v0/z2/z2/z3/temp ;
 wire [3:0] \v0/z2/z2/z4/temp ;
 wire [3:0] \v0/z2/z3/q0 ;
 wire [3:0] \v0/z2/z3/q1 ;
 wire [3:0] \v0/z2/z3/q2 ;
 wire [3:0] \v0/z2/z3/q3 ;
 wire [3:0] \v0/z2/z3/q4 ;
 wire [5:0] \v0/z2/z3/q5 ;
 wire [3:0] \v0/z2/z3/z1/temp ;
 wire [3:0] \v0/z2/z3/z2/temp ;
 wire [3:0] \v0/z2/z3/z3/temp ;
 wire [3:0] \v0/z2/z3/z4/temp ;
 wire [3:0] \v0/z2/z4/q0 ;
 wire [3:0] \v0/z2/z4/q1 ;
 wire [3:0] \v0/z2/z4/q2 ;
 wire [3:0] \v0/z2/z4/q3 ;
 wire [3:0] \v0/z2/z4/q4 ;
 wire [5:0] \v0/z2/z4/q5 ;
 wire [3:0] \v0/z2/z4/z1/temp ;
 wire [3:0] \v0/z2/z4/z2/temp ;
 wire [3:0] \v0/z2/z4/z3/temp ;
 wire [3:0] \v0/z2/z4/z4/temp ;
 wire [7:0] \v0/z3/q0 ;
 wire [7:0] \v0/z3/q1 ;
 wire [7:0] \v0/z3/q2 ;
 wire [7:0] \v0/z3/q3 ;
 wire [7:0] \v0/z3/q4 ;
 wire [11:0] \v0/z3/q5 ;
 wire [3:0] \v0/z3/z1/q0 ;
 wire [3:0] \v0/z3/z1/q1 ;
 wire [3:0] \v0/z3/z1/q2 ;
 wire [3:0] \v0/z3/z1/q3 ;
 wire [3:0] \v0/z3/z1/q4 ;
 wire [5:0] \v0/z3/z1/q5 ;
 wire [3:0] \v0/z3/z1/z1/temp ;
 wire [3:0] \v0/z3/z1/z2/temp ;
 wire [3:0] \v0/z3/z1/z3/temp ;
 wire [3:0] \v0/z3/z1/z4/temp ;
 wire [3:0] \v0/z3/z2/q0 ;
 wire [3:0] \v0/z3/z2/q1 ;
 wire [3:0] \v0/z3/z2/q2 ;
 wire [3:0] \v0/z3/z2/q3 ;
 wire [3:0] \v0/z3/z2/q4 ;
 wire [5:0] \v0/z3/z2/q5 ;
 wire [3:0] \v0/z3/z2/z1/temp ;
 wire [3:0] \v0/z3/z2/z2/temp ;
 wire [3:0] \v0/z3/z2/z3/temp ;
 wire [3:0] \v0/z3/z2/z4/temp ;
 wire [3:0] \v0/z3/z3/q0 ;
 wire [3:0] \v0/z3/z3/q1 ;
 wire [3:0] \v0/z3/z3/q2 ;
 wire [3:0] \v0/z3/z3/q3 ;
 wire [3:0] \v0/z3/z3/q4 ;
 wire [5:0] \v0/z3/z3/q5 ;
 wire [3:0] \v0/z3/z3/z1/temp ;
 wire [3:0] \v0/z3/z3/z2/temp ;
 wire [3:0] \v0/z3/z3/z3/temp ;
 wire [3:0] \v0/z3/z3/z4/temp ;
 wire [3:0] \v0/z3/z4/q0 ;
 wire [3:0] \v0/z3/z4/q1 ;
 wire [3:0] \v0/z3/z4/q2 ;
 wire [3:0] \v0/z3/z4/q3 ;
 wire [3:0] \v0/z3/z4/q4 ;
 wire [5:0] \v0/z3/z4/q5 ;
 wire [3:0] \v0/z3/z4/z1/temp ;
 wire [3:0] \v0/z3/z4/z2/temp ;
 wire [3:0] \v0/z3/z4/z3/temp ;
 wire [3:0] \v0/z3/z4/z4/temp ;
 wire [7:0] \v0/z4/q0 ;
 wire [7:0] \v0/z4/q1 ;
 wire [7:0] \v0/z4/q2 ;
 wire [7:0] \v0/z4/q3 ;
 wire [7:0] \v0/z4/q4 ;
 wire [11:0] \v0/z4/q5 ;
 wire [3:0] \v0/z4/z1/q0 ;
 wire [3:0] \v0/z4/z1/q1 ;
 wire [3:0] \v0/z4/z1/q2 ;
 wire [3:0] \v0/z4/z1/q3 ;
 wire [3:0] \v0/z4/z1/q4 ;
 wire [5:0] \v0/z4/z1/q5 ;
 wire [3:0] \v0/z4/z1/z1/temp ;
 wire [3:0] \v0/z4/z1/z2/temp ;
 wire [3:0] \v0/z4/z1/z3/temp ;
 wire [3:0] \v0/z4/z1/z4/temp ;
 wire [3:0] \v0/z4/z2/q0 ;
 wire [3:0] \v0/z4/z2/q1 ;
 wire [3:0] \v0/z4/z2/q2 ;
 wire [3:0] \v0/z4/z2/q3 ;
 wire [3:0] \v0/z4/z2/q4 ;
 wire [5:0] \v0/z4/z2/q5 ;
 wire [3:0] \v0/z4/z2/z1/temp ;
 wire [3:0] \v0/z4/z2/z2/temp ;
 wire [3:0] \v0/z4/z2/z3/temp ;
 wire [3:0] \v0/z4/z2/z4/temp ;
 wire [3:0] \v0/z4/z3/q0 ;
 wire [3:0] \v0/z4/z3/q1 ;
 wire [3:0] \v0/z4/z3/q2 ;
 wire [3:0] \v0/z4/z3/q3 ;
 wire [3:0] \v0/z4/z3/q4 ;
 wire [5:0] \v0/z4/z3/q5 ;
 wire [3:0] \v0/z4/z3/z1/temp ;
 wire [3:0] \v0/z4/z3/z2/temp ;
 wire [3:0] \v0/z4/z3/z3/temp ;
 wire [3:0] \v0/z4/z3/z4/temp ;
 wire [3:0] \v0/z4/z4/q0 ;
 wire [3:0] \v0/z4/z4/q1 ;
 wire [3:0] \v0/z4/z4/q2 ;
 wire [3:0] \v0/z4/z4/q3 ;
 wire [3:0] \v0/z4/z4/q4 ;
 wire [5:0] \v0/z4/z4/q5 ;
 wire [3:0] \v0/z4/z4/z1/temp ;
 wire [3:0] \v0/z4/z4/z2/temp ;
 wire [3:0] \v0/z4/z4/z3/temp ;
 wire [3:0] \v0/z4/z4/z4/temp ;

 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_65 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_75 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_76 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Left_77 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Right_12 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Left_78 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Right_13 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Left_79 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Right_14 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Left_80 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Right_15 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Left_81 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Right_16 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Left_82 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Right_17 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Left_83 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Right_18 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Left_84 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Right_19 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_66 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Left_85 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Right_20 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Left_86 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Right_21 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Left_87 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Right_22 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Left_88 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Right_23 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Left_89 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Right_24 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Left_90 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Right_25 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Left_91 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Right_26 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Left_92 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Right_27 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Left_93 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Right_28 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Left_94 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Right_29 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_67 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Left_95 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Right_30 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Left_96 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Right_31 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Left_97 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Right_32 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Left_98 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Right_33 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Left_99 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Right_34 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Left_100 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Right_35 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Left_101 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Right_36 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Left_102 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Right_37 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Left_103 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Right_38 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Left_104 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Right_39 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_68 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Left_105 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Right_40 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Left_106 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Right_41 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Left_107 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Right_42 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Left_108 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Right_43 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Left_109 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Right_44 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Left_110 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Right_45 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Left_111 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Right_46 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Left_112 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Right_47 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Left_113 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Right_48 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Left_114 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Right_49 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_69 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Left_115 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Right_50 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Left_116 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Right_51 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Left_117 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Right_52 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Left_118 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Right_53 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Left_119 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Right_54 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Left_120 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Right_55 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Left_121 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Right_56 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Left_122 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Right_57 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Left_123 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Right_58 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Left_124 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Right_59 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_70 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Left_125 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Right_60 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Left_126 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Right_61 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Left_127 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Right_62 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Left_128 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Right_63 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Left_129 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Right_64 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_71 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_72 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_73 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_74 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_228 ();
 sky130_fd_sc_hd__clkinv_1 _072_ (.A(a[1]),
    .Y(_019_));
 sky130_fd_sc_hd__clkinv_1 _073_ (.A(b[1]),
    .Y(_020_));
 sky130_fd_sc_hd__o21ai_0 _074_ (.A1(a[0]),
    .A2(a[1]),
    .B1(a[15]),
    .Y(_021_));
 sky130_fd_sc_hd__a21o_1 _075_ (.A1(a[0]),
    .A2(a[1]),
    .B1(_021_),
    .X(_022_));
 sky130_fd_sc_hd__o21ai_0 _076_ (.A1(_019_),
    .A2(a[15]),
    .B1(_022_),
    .Y(abs_a[1]));
 sky130_fd_sc_hd__xnor2_1 _077_ (.A(a[2]),
    .B(_021_),
    .Y(abs_a[2]));
 sky130_fd_sc_hd__o31ai_1 _078_ (.A1(a[0]),
    .A2(a[1]),
    .A3(a[2]),
    .B1(a[15]),
    .Y(_023_));
 sky130_fd_sc_hd__xnor2_1 _079_ (.A(a[3]),
    .B(_023_),
    .Y(abs_a[3]));
 sky130_fd_sc_hd__or4_1 _080_ (.A(a[0]),
    .B(a[1]),
    .C(a[2]),
    .D(a[3]),
    .X(_024_));
 sky130_fd_sc_hd__nand2_1 _081_ (.A(a[15]),
    .B(_024_),
    .Y(_025_));
 sky130_fd_sc_hd__xnor2_1 _082_ (.A(a[4]),
    .B(_025_),
    .Y(abs_a[4]));
 sky130_fd_sc_hd__o21ai_0 _083_ (.A1(a[4]),
    .A2(_024_),
    .B1(a[15]),
    .Y(_026_));
 sky130_fd_sc_hd__xnor2_1 _084_ (.A(a[5]),
    .B(_026_),
    .Y(abs_a[5]));
 sky130_fd_sc_hd__o31ai_1 _085_ (.A1(a[4]),
    .A2(a[5]),
    .A3(_024_),
    .B1(a[15]),
    .Y(_027_));
 sky130_fd_sc_hd__xnor2_1 _086_ (.A(a[6]),
    .B(_027_),
    .Y(abs_a[6]));
 sky130_fd_sc_hd__nor4_1 _087_ (.A(a[4]),
    .B(a[5]),
    .C(a[6]),
    .D(_024_),
    .Y(_028_));
 sky130_fd_sc_hd__nand2b_1 _088_ (.A_N(_028_),
    .B(a[15]),
    .Y(_029_));
 sky130_fd_sc_hd__xnor2_1 _089_ (.A(a[7]),
    .B(_029_),
    .Y(abs_a[7]));
 sky130_fd_sc_hd__nand2b_1 _090_ (.A_N(a[7]),
    .B(_028_),
    .Y(_030_));
 sky130_fd_sc_hd__nand2_1 _091_ (.A(a[15]),
    .B(_030_),
    .Y(_031_));
 sky130_fd_sc_hd__xnor2_1 _092_ (.A(a[8]),
    .B(_031_),
    .Y(abs_a[8]));
 sky130_fd_sc_hd__o21ai_0 _093_ (.A1(a[8]),
    .A2(_030_),
    .B1(a[15]),
    .Y(_032_));
 sky130_fd_sc_hd__xnor2_1 _094_ (.A(a[9]),
    .B(_032_),
    .Y(abs_a[9]));
 sky130_fd_sc_hd__o31ai_1 _095_ (.A1(a[8]),
    .A2(a[9]),
    .A3(_030_),
    .B1(a[15]),
    .Y(_033_));
 sky130_fd_sc_hd__xnor2_1 _096_ (.A(a[10]),
    .B(_033_),
    .Y(abs_a[10]));
 sky130_fd_sc_hd__or4_1 _097_ (.A(a[8]),
    .B(a[9]),
    .C(a[10]),
    .D(_030_),
    .X(_034_));
 sky130_fd_sc_hd__nand2_1 _098_ (.A(a[15]),
    .B(_034_),
    .Y(_035_));
 sky130_fd_sc_hd__xnor2_1 _099_ (.A(a[11]),
    .B(_035_),
    .Y(abs_a[11]));
 sky130_fd_sc_hd__o21ai_0 _100_ (.A1(a[11]),
    .A2(_034_),
    .B1(a[15]),
    .Y(_036_));
 sky130_fd_sc_hd__xnor2_1 _101_ (.A(a[12]),
    .B(_036_),
    .Y(abs_a[12]));
 sky130_fd_sc_hd__nor3_1 _102_ (.A(a[11]),
    .B(a[12]),
    .C(_034_),
    .Y(_037_));
 sky130_fd_sc_hd__o31ai_1 _103_ (.A1(a[11]),
    .A2(a[12]),
    .A3(_034_),
    .B1(a[15]),
    .Y(_038_));
 sky130_fd_sc_hd__xnor2_1 _104_ (.A(a[13]),
    .B(_038_),
    .Y(abs_a[13]));
 sky130_fd_sc_hd__o41ai_1 _105_ (.A1(a[11]),
    .A2(a[12]),
    .A3(a[13]),
    .A4(_034_),
    .B1(a[15]),
    .Y(_039_));
 sky130_fd_sc_hd__xnor2_1 _106_ (.A(a[14]),
    .B(_039_),
    .Y(abs_a[14]));
 sky130_fd_sc_hd__nor4bb_1 _107_ (.A(a[13]),
    .B(a[14]),
    .C_N(_037_),
    .D_N(a[15]),
    .Y(abs_a[15]));
 sky130_fd_sc_hd__o21ai_0 _108_ (.A1(b[0]),
    .A2(b[1]),
    .B1(b[15]),
    .Y(_000_));
 sky130_fd_sc_hd__a21o_1 _109_ (.A1(b[0]),
    .A2(b[1]),
    .B1(_000_),
    .X(_001_));
 sky130_fd_sc_hd__o21ai_0 _110_ (.A1(_020_),
    .A2(b[15]),
    .B1(_001_),
    .Y(abs_b[1]));
 sky130_fd_sc_hd__xnor2_1 _111_ (.A(b[2]),
    .B(_000_),
    .Y(abs_b[2]));
 sky130_fd_sc_hd__o31ai_1 _112_ (.A1(b[0]),
    .A2(b[1]),
    .A3(b[2]),
    .B1(b[15]),
    .Y(_002_));
 sky130_fd_sc_hd__xnor2_1 _113_ (.A(b[3]),
    .B(_002_),
    .Y(abs_b[3]));
 sky130_fd_sc_hd__or4_1 _114_ (.A(b[0]),
    .B(b[1]),
    .C(b[2]),
    .D(b[3]),
    .X(_003_));
 sky130_fd_sc_hd__nand2_1 _115_ (.A(b[15]),
    .B(_003_),
    .Y(_004_));
 sky130_fd_sc_hd__xnor2_1 _116_ (.A(b[4]),
    .B(_004_),
    .Y(abs_b[4]));
 sky130_fd_sc_hd__o21ai_0 _117_ (.A1(b[4]),
    .A2(_003_),
    .B1(b[15]),
    .Y(_005_));
 sky130_fd_sc_hd__xnor2_1 _118_ (.A(b[5]),
    .B(_005_),
    .Y(abs_b[5]));
 sky130_fd_sc_hd__o31ai_1 _119_ (.A1(b[4]),
    .A2(b[5]),
    .A3(_003_),
    .B1(b[15]),
    .Y(_006_));
 sky130_fd_sc_hd__xnor2_1 _120_ (.A(b[6]),
    .B(_006_),
    .Y(abs_b[6]));
 sky130_fd_sc_hd__nor4_1 _121_ (.A(b[4]),
    .B(b[5]),
    .C(b[6]),
    .D(_003_),
    .Y(_007_));
 sky130_fd_sc_hd__nand2b_1 _122_ (.A_N(_007_),
    .B(b[15]),
    .Y(_008_));
 sky130_fd_sc_hd__xnor2_1 _123_ (.A(b[7]),
    .B(_008_),
    .Y(abs_b[7]));
 sky130_fd_sc_hd__nand2b_1 _124_ (.A_N(b[7]),
    .B(_007_),
    .Y(_009_));
 sky130_fd_sc_hd__nand2_1 _125_ (.A(b[15]),
    .B(_009_),
    .Y(_010_));
 sky130_fd_sc_hd__xnor2_1 _126_ (.A(b[8]),
    .B(_010_),
    .Y(abs_b[8]));
 sky130_fd_sc_hd__o21ai_0 _127_ (.A1(b[8]),
    .A2(_009_),
    .B1(b[15]),
    .Y(_011_));
 sky130_fd_sc_hd__xnor2_1 _128_ (.A(b[9]),
    .B(_011_),
    .Y(abs_b[9]));
 sky130_fd_sc_hd__o31ai_1 _129_ (.A1(b[8]),
    .A2(b[9]),
    .A3(_009_),
    .B1(b[15]),
    .Y(_012_));
 sky130_fd_sc_hd__xnor2_1 _130_ (.A(b[10]),
    .B(_012_),
    .Y(abs_b[10]));
 sky130_fd_sc_hd__or4_1 _131_ (.A(b[8]),
    .B(b[9]),
    .C(b[10]),
    .D(_009_),
    .X(_013_));
 sky130_fd_sc_hd__nand2_1 _132_ (.A(b[15]),
    .B(_013_),
    .Y(_014_));
 sky130_fd_sc_hd__xnor2_1 _133_ (.A(b[11]),
    .B(_014_),
    .Y(abs_b[11]));
 sky130_fd_sc_hd__o21ai_0 _134_ (.A1(b[11]),
    .A2(_013_),
    .B1(b[15]),
    .Y(_015_));
 sky130_fd_sc_hd__xnor2_1 _135_ (.A(b[12]),
    .B(_015_),
    .Y(abs_b[12]));
 sky130_fd_sc_hd__nor3_1 _136_ (.A(b[11]),
    .B(b[12]),
    .C(_013_),
    .Y(_016_));
 sky130_fd_sc_hd__o31ai_1 _137_ (.A1(b[11]),
    .A2(b[12]),
    .A3(_013_),
    .B1(b[15]),
    .Y(_017_));
 sky130_fd_sc_hd__xnor2_1 _138_ (.A(b[13]),
    .B(_017_),
    .Y(abs_b[13]));
 sky130_fd_sc_hd__o41ai_1 _139_ (.A1(b[11]),
    .A2(b[12]),
    .A3(b[13]),
    .A4(_013_),
    .B1(b[15]),
    .Y(_018_));
 sky130_fd_sc_hd__xnor2_1 _140_ (.A(b[14]),
    .B(_018_),
    .Y(abs_b[14]));
 sky130_fd_sc_hd__nor4bb_1 _141_ (.A(b[13]),
    .B(b[14]),
    .C_N(_016_),
    .D_N(b[15]),
    .Y(abs_b[15]));
 sky130_fd_sc_hd__xor2_1 _142_ (.A(a[15]),
    .B(b[15]),
    .X(sign));
 sky130_fd_sc_hd__conb_1 _143_ (.LO(_040_));
 sky130_fd_sc_hd__conb_1 _144_ (.LO(_041_));
 sky130_fd_sc_hd__conb_1 _145_ (.LO(_042_));
 sky130_fd_sc_hd__conb_1 _146_ (.LO(_043_));
 sky130_fd_sc_hd__conb_1 _147_ (.LO(_044_));
 sky130_fd_sc_hd__conb_1 _148_ (.LO(_045_));
 sky130_fd_sc_hd__conb_1 _149_ (.LO(_046_));
 sky130_fd_sc_hd__conb_1 _150_ (.LO(_047_));
 sky130_fd_sc_hd__conb_1 _151_ (.LO(_048_));
 sky130_fd_sc_hd__conb_1 _152_ (.LO(_049_));
 sky130_fd_sc_hd__conb_1 _153_ (.LO(_050_));
 sky130_fd_sc_hd__conb_1 _154_ (.LO(_051_));
 sky130_fd_sc_hd__conb_1 _155_ (.LO(_052_));
 sky130_fd_sc_hd__conb_1 _156_ (.LO(_053_));
 sky130_fd_sc_hd__conb_1 _157_ (.LO(_054_));
 sky130_fd_sc_hd__conb_1 _158_ (.LO(_055_));
 sky130_fd_sc_hd__conb_1 _159_ (.LO(_056_));
 sky130_fd_sc_hd__conb_1 _160_ (.LO(_057_));
 sky130_fd_sc_hd__conb_1 _161_ (.LO(_058_));
 sky130_fd_sc_hd__conb_1 _162_ (.LO(_059_));
 sky130_fd_sc_hd__conb_1 _163_ (.LO(_060_));
 sky130_fd_sc_hd__conb_1 _164_ (.LO(_061_));
 sky130_fd_sc_hd__conb_1 _165_ (.LO(_062_));
 sky130_fd_sc_hd__conb_1 _166_ (.LO(_063_));
 sky130_fd_sc_hd__conb_1 _167_ (.LO(_064_));
 sky130_fd_sc_hd__conb_1 _168_ (.LO(_065_));
 sky130_fd_sc_hd__conb_1 _169_ (.LO(_066_));
 sky130_fd_sc_hd__conb_1 _170_ (.LO(_067_));
 sky130_fd_sc_hd__conb_1 _171_ (.LO(_068_));
 sky130_fd_sc_hd__conb_1 _172_ (.LO(_069_));
 sky130_fd_sc_hd__conb_1 _173_ (.LO(_070_));
 sky130_fd_sc_hd__conb_1 _174_ (.LO(_071_));
 sky130_fd_sc_hd__xor2_1 \inv0/_00_  (.A(sign),
    .B(unsign[0]),
    .X(nextinp[0]));
 sky130_fd_sc_hd__xor2_1 \inv0/_01_  (.A(sign),
    .B(unsign[1]),
    .X(nextinp[1]));
 sky130_fd_sc_hd__xor2_1 \inv0/_02_  (.A(sign),
    .B(unsign[2]),
    .X(nextinp[2]));
 sky130_fd_sc_hd__xor2_1 \inv0/_03_  (.A(sign),
    .B(unsign[3]),
    .X(nextinp[3]));
 sky130_fd_sc_hd__xor2_1 \inv0/_04_  (.A(sign),
    .B(unsign[4]),
    .X(nextinp[4]));
 sky130_fd_sc_hd__xor2_1 \inv0/_05_  (.A(sign),
    .B(unsign[5]),
    .X(nextinp[5]));
 sky130_fd_sc_hd__xor2_1 \inv0/_06_  (.A(sign),
    .B(unsign[6]),
    .X(nextinp[6]));
 sky130_fd_sc_hd__xor2_1 \inv0/_07_  (.A(sign),
    .B(unsign[7]),
    .X(nextinp[7]));
 sky130_fd_sc_hd__xor2_1 \inv0/_08_  (.A(sign),
    .B(unsign[8]),
    .X(nextinp[8]));
 sky130_fd_sc_hd__xor2_1 \inv0/_09_  (.A(sign),
    .B(unsign[9]),
    .X(nextinp[9]));
 sky130_fd_sc_hd__xor2_1 \inv0/_10_  (.A(sign),
    .B(unsign[10]),
    .X(nextinp[10]));
 sky130_fd_sc_hd__xor2_1 \inv0/_11_  (.A(sign),
    .B(unsign[11]),
    .X(nextinp[11]));
 sky130_fd_sc_hd__xor2_1 \inv0/_12_  (.A(sign),
    .B(unsign[12]),
    .X(nextinp[12]));
 sky130_fd_sc_hd__xor2_1 \inv0/_13_  (.A(sign),
    .B(unsign[13]),
    .X(nextinp[13]));
 sky130_fd_sc_hd__xor2_1 \inv0/_14_  (.A(sign),
    .B(unsign[14]),
    .X(nextinp[14]));
 sky130_fd_sc_hd__xor2_1 \inv0/_15_  (.A(sign),
    .B(unsign[15]),
    .X(nextinp[15]));
 sky130_fd_sc_hd__xor2_1 \inv0/_16_  (.A(sign),
    .B(unsign[16]),
    .X(nextinp[16]));
 sky130_fd_sc_hd__xor2_1 \inv0/_17_  (.A(sign),
    .B(unsign[17]),
    .X(nextinp[17]));
 sky130_fd_sc_hd__xor2_1 \inv0/_18_  (.A(sign),
    .B(unsign[18]),
    .X(nextinp[18]));
 sky130_fd_sc_hd__xor2_1 \inv0/_19_  (.A(sign),
    .B(unsign[19]),
    .X(nextinp[19]));
 sky130_fd_sc_hd__xor2_1 \inv0/_20_  (.A(sign),
    .B(unsign[20]),
    .X(nextinp[20]));
 sky130_fd_sc_hd__xor2_1 \inv0/_21_  (.A(sign),
    .B(unsign[21]),
    .X(nextinp[21]));
 sky130_fd_sc_hd__xor2_1 \inv0/_22_  (.A(sign),
    .B(unsign[22]),
    .X(nextinp[22]));
 sky130_fd_sc_hd__xor2_1 \inv0/_23_  (.A(sign),
    .B(unsign[23]),
    .X(nextinp[23]));
 sky130_fd_sc_hd__xor2_1 \inv0/_24_  (.A(sign),
    .B(unsign[24]),
    .X(nextinp[24]));
 sky130_fd_sc_hd__xor2_1 \inv0/_25_  (.A(sign),
    .B(unsign[25]),
    .X(nextinp[25]));
 sky130_fd_sc_hd__xor2_1 \inv0/_26_  (.A(sign),
    .B(unsign[26]),
    .X(nextinp[26]));
 sky130_fd_sc_hd__xor2_1 \inv0/_27_  (.A(sign),
    .B(unsign[27]),
    .X(nextinp[27]));
 sky130_fd_sc_hd__xor2_1 \inv0/_28_  (.A(sign),
    .B(unsign[28]),
    .X(nextinp[28]));
 sky130_fd_sc_hd__xor2_1 \inv0/_29_  (.A(sign),
    .B(unsign[29]),
    .X(nextinp[29]));
 sky130_fd_sc_hd__xor2_1 \inv0/_30_  (.A(sign),
    .B(unsign[30]),
    .X(nextinp[30]));
 sky130_fd_sc_hd__xor2_1 \inv0/_31_  (.A(sign),
    .B(unsign[31]),
    .X(nextinp[31]));
 sky130_fd_sc_hd__xnor2_1 \lastadder/ksa32/_163_  (.A(_040_),
    .B(nextinp[0]),
    .Y(\lastadder/ksa32/_162_ ));
 sky130_fd_sc_hd__xnor2_1 \lastadder/ksa32/_164_  (.A(sign),
    .B(\lastadder/ksa32/_162_ ),
    .Y(c[0]));
 sky130_fd_sc_hd__maj3_1 \lastadder/ksa32/_165_  (.A(_040_),
    .B(nextinp[0]),
    .C(sign),
    .X(\lastadder/ksa32/_000_ ));
 sky130_fd_sc_hd__lpflow_inputiso1p_1 \lastadder/ksa32/_166_  (.A(_041_),
    .SLEEP(nextinp[1]),
    .X(\lastadder/ksa32/_001_ ));
 sky130_fd_sc_hd__and2_0 \lastadder/ksa32/_167_  (.A(_041_),
    .B(nextinp[1]),
    .X(\lastadder/ksa32/_002_ ));
 sky130_fd_sc_hd__nand2_1 \lastadder/ksa32/_168_  (.A(_041_),
    .B(nextinp[1]),
    .Y(\lastadder/ksa32/_003_ ));
 sky130_fd_sc_hd__nand2_1 \lastadder/ksa32/_169_  (.A(\lastadder/ksa32/_001_ ),
    .B(\lastadder/ksa32/_003_ ),
    .Y(\lastadder/ksa32/_004_ ));
 sky130_fd_sc_hd__xnor2_1 \lastadder/ksa32/_170_  (.A(\lastadder/ksa32/_000_ ),
    .B(\lastadder/ksa32/_004_ ),
    .Y(c[1]));
 sky130_fd_sc_hd__nor2_1 \lastadder/ksa32/_171_  (.A(_042_),
    .B(nextinp[2]),
    .Y(\lastadder/ksa32/_005_ ));
 sky130_fd_sc_hd__xor2_1 \lastadder/ksa32/_172_  (.A(_042_),
    .B(nextinp[2]),
    .X(\lastadder/ksa32/_006_ ));
 sky130_fd_sc_hd__a21oi_1 \lastadder/ksa32/_173_  (.A1(\lastadder/ksa32/_000_ ),
    .A2(\lastadder/ksa32/_001_ ),
    .B1(\lastadder/ksa32/_002_ ),
    .Y(\lastadder/ksa32/_007_ ));
 sky130_fd_sc_hd__xnor2_1 \lastadder/ksa32/_174_  (.A(\lastadder/ksa32/_006_ ),
    .B(\lastadder/ksa32/_007_ ),
    .Y(c[2]));
 sky130_fd_sc_hd__nand2_1 \lastadder/ksa32/_175_  (.A(_043_),
    .B(nextinp[3]),
    .Y(\lastadder/ksa32/_008_ ));
 sky130_fd_sc_hd__xnor2_1 \lastadder/ksa32/_176_  (.A(_043_),
    .B(nextinp[3]),
    .Y(\lastadder/ksa32/_009_ ));
 sky130_fd_sc_hd__a221oi_1 \lastadder/ksa32/_177_  (.A1(_042_),
    .A2(nextinp[2]),
    .B1(\lastadder/ksa32/_000_ ),
    .B2(\lastadder/ksa32/_001_ ),
    .C1(\lastadder/ksa32/_002_ ),
    .Y(\lastadder/ksa32/_010_ ));
 sky130_fd_sc_hd__o21a_1 \lastadder/ksa32/_178_  (.A1(\lastadder/ksa32/_005_ ),
    .A2(\lastadder/ksa32/_010_ ),
    .B1(\lastadder/ksa32/_009_ ),
    .X(\lastadder/ksa32/_011_ ));
 sky130_fd_sc_hd__nor3_1 \lastadder/ksa32/_179_  (.A(\lastadder/ksa32/_005_ ),
    .B(\lastadder/ksa32/_009_ ),
    .C(\lastadder/ksa32/_010_ ),
    .Y(\lastadder/ksa32/_012_ ));
 sky130_fd_sc_hd__nor2_1 \lastadder/ksa32/_180_  (.A(\lastadder/ksa32/_011_ ),
    .B(\lastadder/ksa32/_012_ ),
    .Y(c[3]));
 sky130_fd_sc_hd__lpflow_inputiso1p_1 \lastadder/ksa32/_181_  (.A(_044_),
    .SLEEP(nextinp[4]),
    .X(\lastadder/ksa32/_013_ ));
 sky130_fd_sc_hd__nand2_1 \lastadder/ksa32/_182_  (.A(_044_),
    .B(nextinp[4]),
    .Y(\lastadder/ksa32/_014_ ));
 sky130_fd_sc_hd__nand2_1 \lastadder/ksa32/_183_  (.A(\lastadder/ksa32/_013_ ),
    .B(\lastadder/ksa32/_014_ ),
    .Y(\lastadder/ksa32/_015_ ));
 sky130_fd_sc_hd__a21oi_1 \lastadder/ksa32/_184_  (.A1(_043_),
    .A2(nextinp[3]),
    .B1(\lastadder/ksa32/_012_ ),
    .Y(\lastadder/ksa32/_016_ ));
 sky130_fd_sc_hd__xor2_1 \lastadder/ksa32/_185_  (.A(\lastadder/ksa32/_015_ ),
    .B(\lastadder/ksa32/_016_ ),
    .X(c[4]));
 sky130_fd_sc_hd__lpflow_inputiso1p_1 \lastadder/ksa32/_186_  (.A(_045_),
    .SLEEP(nextinp[5]),
    .X(\lastadder/ksa32/_017_ ));
 sky130_fd_sc_hd__and2_0 \lastadder/ksa32/_187_  (.A(_045_),
    .B(nextinp[5]),
    .X(\lastadder/ksa32/_018_ ));
 sky130_fd_sc_hd__nand2_1 \lastadder/ksa32/_188_  (.A(_045_),
    .B(nextinp[5]),
    .Y(\lastadder/ksa32/_019_ ));
 sky130_fd_sc_hd__nand2_1 \lastadder/ksa32/_189_  (.A(\lastadder/ksa32/_017_ ),
    .B(\lastadder/ksa32/_019_ ),
    .Y(\lastadder/ksa32/_020_ ));
 sky130_fd_sc_hd__o311ai_0 \lastadder/ksa32/_190_  (.A1(\lastadder/ksa32/_005_ ),
    .A2(\lastadder/ksa32/_009_ ),
    .A3(\lastadder/ksa32/_010_ ),
    .B1(\lastadder/ksa32/_014_ ),
    .C1(\lastadder/ksa32/_008_ ),
    .Y(\lastadder/ksa32/_021_ ));
 sky130_fd_sc_hd__and2_0 \lastadder/ksa32/_191_  (.A(\lastadder/ksa32/_013_ ),
    .B(\lastadder/ksa32/_021_ ),
    .X(\lastadder/ksa32/_022_ ));
 sky130_fd_sc_hd__xnor2_1 \lastadder/ksa32/_192_  (.A(\lastadder/ksa32/_020_ ),
    .B(\lastadder/ksa32/_022_ ),
    .Y(c[5]));
 sky130_fd_sc_hd__a21oi_1 \lastadder/ksa32/_193_  (.A1(\lastadder/ksa32/_017_ ),
    .A2(\lastadder/ksa32/_022_ ),
    .B1(\lastadder/ksa32/_018_ ),
    .Y(\lastadder/ksa32/_023_ ));
 sky130_fd_sc_hd__nor2_1 \lastadder/ksa32/_194_  (.A(_046_),
    .B(nextinp[6]),
    .Y(\lastadder/ksa32/_024_ ));
 sky130_fd_sc_hd__and2_0 \lastadder/ksa32/_195_  (.A(_046_),
    .B(nextinp[6]),
    .X(\lastadder/ksa32/_025_ ));
 sky130_fd_sc_hd__nor2_1 \lastadder/ksa32/_196_  (.A(\lastadder/ksa32/_024_ ),
    .B(\lastadder/ksa32/_025_ ),
    .Y(\lastadder/ksa32/_026_ ));
 sky130_fd_sc_hd__xnor2_1 \lastadder/ksa32/_197_  (.A(\lastadder/ksa32/_023_ ),
    .B(\lastadder/ksa32/_026_ ),
    .Y(c[6]));
 sky130_fd_sc_hd__nor2_1 \lastadder/ksa32/_198_  (.A(_047_),
    .B(nextinp[7]),
    .Y(\lastadder/ksa32/_027_ ));
 sky130_fd_sc_hd__nand2_1 \lastadder/ksa32/_199_  (.A(_047_),
    .B(nextinp[7]),
    .Y(\lastadder/ksa32/_028_ ));
 sky130_fd_sc_hd__nand2b_1 \lastadder/ksa32/_200_  (.A_N(\lastadder/ksa32/_027_ ),
    .B(\lastadder/ksa32/_028_ ),
    .Y(\lastadder/ksa32/_029_ ));
 sky130_fd_sc_hd__a311oi_1 \lastadder/ksa32/_201_  (.A1(\lastadder/ksa32/_013_ ),
    .A2(\lastadder/ksa32/_017_ ),
    .A3(\lastadder/ksa32/_021_ ),
    .B1(\lastadder/ksa32/_025_ ),
    .C1(\lastadder/ksa32/_018_ ),
    .Y(\lastadder/ksa32/_030_ ));
 sky130_fd_sc_hd__nor2_1 \lastadder/ksa32/_202_  (.A(\lastadder/ksa32/_024_ ),
    .B(\lastadder/ksa32/_030_ ),
    .Y(\lastadder/ksa32/_031_ ));
 sky130_fd_sc_hd__xnor2_1 \lastadder/ksa32/_203_  (.A(\lastadder/ksa32/_029_ ),
    .B(\lastadder/ksa32/_031_ ),
    .Y(c[7]));
 sky130_fd_sc_hd__nor2_1 \lastadder/ksa32/_204_  (.A(_048_),
    .B(nextinp[8]),
    .Y(\lastadder/ksa32/_032_ ));
 sky130_fd_sc_hd__and2_0 \lastadder/ksa32/_205_  (.A(_048_),
    .B(nextinp[8]),
    .X(\lastadder/ksa32/_033_ ));
 sky130_fd_sc_hd__nand2_1 \lastadder/ksa32/_206_  (.A(_048_),
    .B(nextinp[8]),
    .Y(\lastadder/ksa32/_034_ ));
 sky130_fd_sc_hd__o31a_1 \lastadder/ksa32/_207_  (.A1(\lastadder/ksa32/_024_ ),
    .A2(\lastadder/ksa32/_027_ ),
    .A3(\lastadder/ksa32/_030_ ),
    .B1(\lastadder/ksa32/_028_ ),
    .X(\lastadder/ksa32/_035_ ));
 sky130_fd_sc_hd__or3_1 \lastadder/ksa32/_208_  (.A(\lastadder/ksa32/_032_ ),
    .B(\lastadder/ksa32/_033_ ),
    .C(\lastadder/ksa32/_035_ ),
    .X(\lastadder/ksa32/_036_ ));
 sky130_fd_sc_hd__o21ai_0 \lastadder/ksa32/_209_  (.A1(\lastadder/ksa32/_032_ ),
    .A2(\lastadder/ksa32/_033_ ),
    .B1(\lastadder/ksa32/_035_ ),
    .Y(\lastadder/ksa32/_037_ ));
 sky130_fd_sc_hd__and2_0 \lastadder/ksa32/_210_  (.A(\lastadder/ksa32/_036_ ),
    .B(\lastadder/ksa32/_037_ ),
    .X(c[8]));
 sky130_fd_sc_hd__nor2_1 \lastadder/ksa32/_211_  (.A(_049_),
    .B(nextinp[9]),
    .Y(\lastadder/ksa32/_038_ ));
 sky130_fd_sc_hd__nand2_1 \lastadder/ksa32/_212_  (.A(_049_),
    .B(nextinp[9]),
    .Y(\lastadder/ksa32/_039_ ));
 sky130_fd_sc_hd__nor2b_1 \lastadder/ksa32/_213_  (.A(\lastadder/ksa32/_038_ ),
    .B_N(\lastadder/ksa32/_039_ ),
    .Y(\lastadder/ksa32/_040_ ));
 sky130_fd_sc_hd__o311a_1 \lastadder/ksa32/_214_  (.A1(\lastadder/ksa32/_024_ ),
    .A2(\lastadder/ksa32/_027_ ),
    .A3(\lastadder/ksa32/_030_ ),
    .B1(\lastadder/ksa32/_034_ ),
    .C1(\lastadder/ksa32/_028_ ),
    .X(\lastadder/ksa32/_041_ ));
 sky130_fd_sc_hd__nor2_1 \lastadder/ksa32/_215_  (.A(\lastadder/ksa32/_032_ ),
    .B(\lastadder/ksa32/_041_ ),
    .Y(\lastadder/ksa32/_042_ ));
 sky130_fd_sc_hd__xor2_1 \lastadder/ksa32/_216_  (.A(\lastadder/ksa32/_040_ ),
    .B(\lastadder/ksa32/_042_ ),
    .X(c[9]));
 sky130_fd_sc_hd__nor2_1 \lastadder/ksa32/_217_  (.A(_050_),
    .B(nextinp[10]),
    .Y(\lastadder/ksa32/_043_ ));
 sky130_fd_sc_hd__nand2_1 \lastadder/ksa32/_218_  (.A(_050_),
    .B(nextinp[10]),
    .Y(\lastadder/ksa32/_044_ ));
 sky130_fd_sc_hd__nand2b_1 \lastadder/ksa32/_219_  (.A_N(\lastadder/ksa32/_043_ ),
    .B(\lastadder/ksa32/_044_ ),
    .Y(\lastadder/ksa32/_045_ ));
 sky130_fd_sc_hd__a31oi_1 \lastadder/ksa32/_220_  (.A1(\lastadder/ksa32/_034_ ),
    .A2(\lastadder/ksa32/_036_ ),
    .A3(\lastadder/ksa32/_039_ ),
    .B1(\lastadder/ksa32/_038_ ),
    .Y(\lastadder/ksa32/_046_ ));
 sky130_fd_sc_hd__nand2b_1 \lastadder/ksa32/_221_  (.A_N(\lastadder/ksa32/_045_ ),
    .B(\lastadder/ksa32/_046_ ),
    .Y(\lastadder/ksa32/_047_ ));
 sky130_fd_sc_hd__xnor2_1 \lastadder/ksa32/_222_  (.A(\lastadder/ksa32/_045_ ),
    .B(\lastadder/ksa32/_046_ ),
    .Y(c[10]));
 sky130_fd_sc_hd__nor2_1 \lastadder/ksa32/_223_  (.A(_051_),
    .B(nextinp[11]),
    .Y(\lastadder/ksa32/_048_ ));
 sky130_fd_sc_hd__nand2_1 \lastadder/ksa32/_224_  (.A(_051_),
    .B(nextinp[11]),
    .Y(\lastadder/ksa32/_049_ ));
 sky130_fd_sc_hd__nand2b_1 \lastadder/ksa32/_225_  (.A_N(\lastadder/ksa32/_048_ ),
    .B(\lastadder/ksa32/_049_ ),
    .Y(\lastadder/ksa32/_050_ ));
 sky130_fd_sc_hd__o311a_1 \lastadder/ksa32/_226_  (.A1(\lastadder/ksa32/_032_ ),
    .A2(\lastadder/ksa32/_038_ ),
    .A3(\lastadder/ksa32/_041_ ),
    .B1(\lastadder/ksa32/_044_ ),
    .C1(\lastadder/ksa32/_039_ ),
    .X(\lastadder/ksa32/_051_ ));
 sky130_fd_sc_hd__nor2_1 \lastadder/ksa32/_227_  (.A(\lastadder/ksa32/_043_ ),
    .B(\lastadder/ksa32/_051_ ),
    .Y(\lastadder/ksa32/_052_ ));
 sky130_fd_sc_hd__xnor2_1 \lastadder/ksa32/_228_  (.A(\lastadder/ksa32/_050_ ),
    .B(\lastadder/ksa32/_052_ ),
    .Y(c[11]));
 sky130_fd_sc_hd__nor2_1 \lastadder/ksa32/_229_  (.A(_052_),
    .B(nextinp[12]),
    .Y(\lastadder/ksa32/_053_ ));
 sky130_fd_sc_hd__nand2_1 \lastadder/ksa32/_230_  (.A(_052_),
    .B(nextinp[12]),
    .Y(\lastadder/ksa32/_054_ ));
 sky130_fd_sc_hd__nor2b_1 \lastadder/ksa32/_231_  (.A(\lastadder/ksa32/_053_ ),
    .B_N(\lastadder/ksa32/_054_ ),
    .Y(\lastadder/ksa32/_055_ ));
 sky130_fd_sc_hd__clkinv_1 \lastadder/ksa32/_232_  (.A(\lastadder/ksa32/_055_ ),
    .Y(\lastadder/ksa32/_056_ ));
 sky130_fd_sc_hd__a31oi_1 \lastadder/ksa32/_233_  (.A1(\lastadder/ksa32/_044_ ),
    .A2(\lastadder/ksa32/_047_ ),
    .A3(\lastadder/ksa32/_049_ ),
    .B1(\lastadder/ksa32/_048_ ),
    .Y(\lastadder/ksa32/_057_ ));
 sky130_fd_sc_hd__xnor2_1 \lastadder/ksa32/_234_  (.A(\lastadder/ksa32/_056_ ),
    .B(\lastadder/ksa32/_057_ ),
    .Y(c[12]));
 sky130_fd_sc_hd__nor2_1 \lastadder/ksa32/_235_  (.A(_053_),
    .B(nextinp[13]),
    .Y(\lastadder/ksa32/_058_ ));
 sky130_fd_sc_hd__nand2_1 \lastadder/ksa32/_236_  (.A(_053_),
    .B(nextinp[13]),
    .Y(\lastadder/ksa32/_059_ ));
 sky130_fd_sc_hd__nor2b_1 \lastadder/ksa32/_237_  (.A(\lastadder/ksa32/_058_ ),
    .B_N(\lastadder/ksa32/_059_ ),
    .Y(\lastadder/ksa32/_060_ ));
 sky130_fd_sc_hd__a21o_1 \lastadder/ksa32/_238_  (.A1(\lastadder/ksa32/_049_ ),
    .A2(\lastadder/ksa32/_054_ ),
    .B1(\lastadder/ksa32/_053_ ),
    .X(\lastadder/ksa32/_061_ ));
 sky130_fd_sc_hd__o41ai_1 \lastadder/ksa32/_239_  (.A1(\lastadder/ksa32/_043_ ),
    .A2(\lastadder/ksa32/_050_ ),
    .A3(\lastadder/ksa32/_051_ ),
    .A4(\lastadder/ksa32/_056_ ),
    .B1(\lastadder/ksa32/_061_ ),
    .Y(\lastadder/ksa32/_062_ ));
 sky130_fd_sc_hd__xor2_1 \lastadder/ksa32/_240_  (.A(\lastadder/ksa32/_060_ ),
    .B(\lastadder/ksa32/_062_ ),
    .X(c[13]));
 sky130_fd_sc_hd__nor2_1 \lastadder/ksa32/_241_  (.A(_054_),
    .B(nextinp[14]),
    .Y(\lastadder/ksa32/_063_ ));
 sky130_fd_sc_hd__nand2_1 \lastadder/ksa32/_242_  (.A(_054_),
    .B(nextinp[14]),
    .Y(\lastadder/ksa32/_064_ ));
 sky130_fd_sc_hd__nor2b_1 \lastadder/ksa32/_243_  (.A(\lastadder/ksa32/_063_ ),
    .B_N(\lastadder/ksa32/_064_ ),
    .Y(\lastadder/ksa32/_065_ ));
 sky130_fd_sc_hd__o21ai_0 \lastadder/ksa32/_244_  (.A1(\lastadder/ksa32/_054_ ),
    .A2(\lastadder/ksa32/_058_ ),
    .B1(\lastadder/ksa32/_059_ ),
    .Y(\lastadder/ksa32/_066_ ));
 sky130_fd_sc_hd__a31oi_1 \lastadder/ksa32/_245_  (.A1(\lastadder/ksa32/_055_ ),
    .A2(\lastadder/ksa32/_057_ ),
    .A3(\lastadder/ksa32/_060_ ),
    .B1(\lastadder/ksa32/_066_ ),
    .Y(\lastadder/ksa32/_067_ ));
 sky130_fd_sc_hd__xnor2_1 \lastadder/ksa32/_246_  (.A(\lastadder/ksa32/_065_ ),
    .B(\lastadder/ksa32/_067_ ),
    .Y(c[14]));
 sky130_fd_sc_hd__nor2_1 \lastadder/ksa32/_247_  (.A(_055_),
    .B(nextinp[15]),
    .Y(\lastadder/ksa32/_068_ ));
 sky130_fd_sc_hd__nand2_1 \lastadder/ksa32/_248_  (.A(_055_),
    .B(nextinp[15]),
    .Y(\lastadder/ksa32/_069_ ));
 sky130_fd_sc_hd__nor2b_1 \lastadder/ksa32/_249_  (.A(\lastadder/ksa32/_068_ ),
    .B_N(\lastadder/ksa32/_069_ ),
    .Y(\lastadder/ksa32/_070_ ));
 sky130_fd_sc_hd__a21oi_1 \lastadder/ksa32/_250_  (.A1(\lastadder/ksa32/_059_ ),
    .A2(\lastadder/ksa32/_064_ ),
    .B1(\lastadder/ksa32/_063_ ),
    .Y(\lastadder/ksa32/_071_ ));
 sky130_fd_sc_hd__a31oi_1 \lastadder/ksa32/_251_  (.A1(\lastadder/ksa32/_060_ ),
    .A2(\lastadder/ksa32/_062_ ),
    .A3(\lastadder/ksa32/_065_ ),
    .B1(\lastadder/ksa32/_071_ ),
    .Y(\lastadder/ksa32/_072_ ));
 sky130_fd_sc_hd__xnor2_1 \lastadder/ksa32/_252_  (.A(\lastadder/ksa32/_070_ ),
    .B(\lastadder/ksa32/_072_ ),
    .Y(c[15]));
 sky130_fd_sc_hd__nor2_1 \lastadder/ksa32/_253_  (.A(_056_),
    .B(nextinp[16]),
    .Y(\lastadder/ksa32/_073_ ));
 sky130_fd_sc_hd__nand2_1 \lastadder/ksa32/_254_  (.A(_056_),
    .B(nextinp[16]),
    .Y(\lastadder/ksa32/_074_ ));
 sky130_fd_sc_hd__nor2b_1 \lastadder/ksa32/_255_  (.A(\lastadder/ksa32/_073_ ),
    .B_N(\lastadder/ksa32/_074_ ),
    .Y(\lastadder/ksa32/_075_ ));
 sky130_fd_sc_hd__o211ai_1 \lastadder/ksa32/_256_  (.A1(\lastadder/ksa32/_063_ ),
    .A2(\lastadder/ksa32/_067_ ),
    .B1(\lastadder/ksa32/_069_ ),
    .C1(\lastadder/ksa32/_064_ ),
    .Y(\lastadder/ksa32/_076_ ));
 sky130_fd_sc_hd__o21ai_0 \lastadder/ksa32/_257_  (.A1(_055_),
    .A2(nextinp[15]),
    .B1(\lastadder/ksa32/_076_ ),
    .Y(\lastadder/ksa32/_077_ ));
 sky130_fd_sc_hd__xnor2_1 \lastadder/ksa32/_258_  (.A(\lastadder/ksa32/_075_ ),
    .B(\lastadder/ksa32/_077_ ),
    .Y(c[16]));
 sky130_fd_sc_hd__nand2_1 \lastadder/ksa32/_259_  (.A(_057_),
    .B(nextinp[17]),
    .Y(\lastadder/ksa32/_078_ ));
 sky130_fd_sc_hd__xnor2_1 \lastadder/ksa32/_260_  (.A(_057_),
    .B(nextinp[17]),
    .Y(\lastadder/ksa32/_079_ ));
 sky130_fd_sc_hd__o211a_1 \lastadder/ksa32/_261_  (.A1(\lastadder/ksa32/_068_ ),
    .A2(\lastadder/ksa32/_072_ ),
    .B1(\lastadder/ksa32/_074_ ),
    .C1(\lastadder/ksa32/_069_ ),
    .X(\lastadder/ksa32/_080_ ));
 sky130_fd_sc_hd__nor2_1 \lastadder/ksa32/_262_  (.A(\lastadder/ksa32/_073_ ),
    .B(\lastadder/ksa32/_080_ ),
    .Y(\lastadder/ksa32/_081_ ));
 sky130_fd_sc_hd__nor3_1 \lastadder/ksa32/_263_  (.A(\lastadder/ksa32/_073_ ),
    .B(\lastadder/ksa32/_079_ ),
    .C(\lastadder/ksa32/_080_ ),
    .Y(\lastadder/ksa32/_082_ ));
 sky130_fd_sc_hd__xnor2_1 \lastadder/ksa32/_264_  (.A(\lastadder/ksa32/_079_ ),
    .B(\lastadder/ksa32/_081_ ),
    .Y(c[17]));
 sky130_fd_sc_hd__nor2_1 \lastadder/ksa32/_265_  (.A(_058_),
    .B(nextinp[18]),
    .Y(\lastadder/ksa32/_083_ ));
 sky130_fd_sc_hd__nand2_1 \lastadder/ksa32/_266_  (.A(_058_),
    .B(nextinp[18]),
    .Y(\lastadder/ksa32/_084_ ));
 sky130_fd_sc_hd__nor2b_1 \lastadder/ksa32/_267_  (.A(\lastadder/ksa32/_083_ ),
    .B_N(\lastadder/ksa32/_084_ ),
    .Y(\lastadder/ksa32/_085_ ));
 sky130_fd_sc_hd__o31a_1 \lastadder/ksa32/_268_  (.A1(\lastadder/ksa32/_073_ ),
    .A2(\lastadder/ksa32/_079_ ),
    .A3(\lastadder/ksa32/_080_ ),
    .B1(\lastadder/ksa32/_078_ ),
    .X(\lastadder/ksa32/_086_ ));
 sky130_fd_sc_hd__xnor2_1 \lastadder/ksa32/_269_  (.A(\lastadder/ksa32/_085_ ),
    .B(\lastadder/ksa32/_086_ ),
    .Y(c[18]));
 sky130_fd_sc_hd__nor2_1 \lastadder/ksa32/_270_  (.A(_059_),
    .B(nextinp[19]),
    .Y(\lastadder/ksa32/_087_ ));
 sky130_fd_sc_hd__xor2_1 \lastadder/ksa32/_271_  (.A(_059_),
    .B(nextinp[19]),
    .X(\lastadder/ksa32/_088_ ));
 sky130_fd_sc_hd__nand2_1 \lastadder/ksa32/_272_  (.A(\lastadder/ksa32/_078_ ),
    .B(\lastadder/ksa32/_084_ ),
    .Y(\lastadder/ksa32/_089_ ));
 sky130_fd_sc_hd__o21ai_0 \lastadder/ksa32/_273_  (.A1(\lastadder/ksa32/_083_ ),
    .A2(\lastadder/ksa32/_086_ ),
    .B1(\lastadder/ksa32/_084_ ),
    .Y(\lastadder/ksa32/_090_ ));
 sky130_fd_sc_hd__o221ai_1 \lastadder/ksa32/_274_  (.A1(_058_),
    .A2(nextinp[18]),
    .B1(\lastadder/ksa32/_082_ ),
    .B2(\lastadder/ksa32/_089_ ),
    .C1(\lastadder/ksa32/_088_ ),
    .Y(\lastadder/ksa32/_091_ ));
 sky130_fd_sc_hd__xor2_1 \lastadder/ksa32/_275_  (.A(\lastadder/ksa32/_088_ ),
    .B(\lastadder/ksa32/_090_ ),
    .X(c[19]));
 sky130_fd_sc_hd__nor2_1 \lastadder/ksa32/_276_  (.A(_060_),
    .B(nextinp[20]),
    .Y(\lastadder/ksa32/_092_ ));
 sky130_fd_sc_hd__nand2_1 \lastadder/ksa32/_277_  (.A(_060_),
    .B(nextinp[20]),
    .Y(\lastadder/ksa32/_093_ ));
 sky130_fd_sc_hd__nand2b_1 \lastadder/ksa32/_278_  (.A_N(\lastadder/ksa32/_092_ ),
    .B(\lastadder/ksa32/_093_ ),
    .Y(\lastadder/ksa32/_094_ ));
 sky130_fd_sc_hd__clkinv_1 \lastadder/ksa32/_279_  (.A(\lastadder/ksa32/_094_ ),
    .Y(\lastadder/ksa32/_095_ ));
 sky130_fd_sc_hd__nand2_1 \lastadder/ksa32/_280_  (.A(\lastadder/ksa32/_085_ ),
    .B(\lastadder/ksa32/_088_ ),
    .Y(\lastadder/ksa32/_096_ ));
 sky130_fd_sc_hd__nor2_1 \lastadder/ksa32/_281_  (.A(\lastadder/ksa32/_084_ ),
    .B(\lastadder/ksa32/_087_ ),
    .Y(\lastadder/ksa32/_097_ ));
 sky130_fd_sc_hd__a21oi_1 \lastadder/ksa32/_282_  (.A1(_059_),
    .A2(nextinp[19]),
    .B1(\lastadder/ksa32/_097_ ),
    .Y(\lastadder/ksa32/_098_ ));
 sky130_fd_sc_hd__o21ai_0 \lastadder/ksa32/_283_  (.A1(\lastadder/ksa32/_086_ ),
    .A2(\lastadder/ksa32/_096_ ),
    .B1(\lastadder/ksa32/_098_ ),
    .Y(\lastadder/ksa32/_099_ ));
 sky130_fd_sc_hd__xnor2_1 \lastadder/ksa32/_284_  (.A(\lastadder/ksa32/_094_ ),
    .B(\lastadder/ksa32/_099_ ),
    .Y(c[20]));
 sky130_fd_sc_hd__nor2_1 \lastadder/ksa32/_285_  (.A(_061_),
    .B(nextinp[21]),
    .Y(\lastadder/ksa32/_100_ ));
 sky130_fd_sc_hd__nand2_1 \lastadder/ksa32/_286_  (.A(_061_),
    .B(nextinp[21]),
    .Y(\lastadder/ksa32/_101_ ));
 sky130_fd_sc_hd__nor2b_1 \lastadder/ksa32/_287_  (.A(\lastadder/ksa32/_100_ ),
    .B_N(\lastadder/ksa32/_101_ ),
    .Y(\lastadder/ksa32/_102_ ));
 sky130_fd_sc_hd__clkinv_1 \lastadder/ksa32/_288_  (.A(\lastadder/ksa32/_102_ ),
    .Y(\lastadder/ksa32/_103_ ));
 sky130_fd_sc_hd__a22oi_1 \lastadder/ksa32/_289_  (.A1(_059_),
    .A2(nextinp[19]),
    .B1(_060_),
    .B2(nextinp[20]),
    .Y(\lastadder/ksa32/_104_ ));
 sky130_fd_sc_hd__a21oi_1 \lastadder/ksa32/_290_  (.A1(\lastadder/ksa32/_091_ ),
    .A2(\lastadder/ksa32/_104_ ),
    .B1(\lastadder/ksa32/_092_ ),
    .Y(\lastadder/ksa32/_105_ ));
 sky130_fd_sc_hd__nor2_1 \lastadder/ksa32/_291_  (.A(\lastadder/ksa32/_102_ ),
    .B(\lastadder/ksa32/_105_ ),
    .Y(\lastadder/ksa32/_106_ ));
 sky130_fd_sc_hd__a211oi_1 \lastadder/ksa32/_292_  (.A1(\lastadder/ksa32/_091_ ),
    .A2(\lastadder/ksa32/_104_ ),
    .B1(\lastadder/ksa32/_103_ ),
    .C1(\lastadder/ksa32/_092_ ),
    .Y(\lastadder/ksa32/_107_ ));
 sky130_fd_sc_hd__nor2_1 \lastadder/ksa32/_293_  (.A(\lastadder/ksa32/_106_ ),
    .B(\lastadder/ksa32/_107_ ),
    .Y(c[21]));
 sky130_fd_sc_hd__lpflow_inputiso1p_1 \lastadder/ksa32/_294_  (.A(_062_),
    .SLEEP(nextinp[22]),
    .X(\lastadder/ksa32/_108_ ));
 sky130_fd_sc_hd__nand2_1 \lastadder/ksa32/_295_  (.A(_062_),
    .B(nextinp[22]),
    .Y(\lastadder/ksa32/_109_ ));
 sky130_fd_sc_hd__and2_0 \lastadder/ksa32/_296_  (.A(\lastadder/ksa32/_108_ ),
    .B(\lastadder/ksa32/_109_ ),
    .X(\lastadder/ksa32/_110_ ));
 sky130_fd_sc_hd__o21ai_0 \lastadder/ksa32/_297_  (.A1(\lastadder/ksa32/_093_ ),
    .A2(\lastadder/ksa32/_100_ ),
    .B1(\lastadder/ksa32/_101_ ),
    .Y(\lastadder/ksa32/_111_ ));
 sky130_fd_sc_hd__a31oi_1 \lastadder/ksa32/_298_  (.A1(\lastadder/ksa32/_095_ ),
    .A2(\lastadder/ksa32/_099_ ),
    .A3(\lastadder/ksa32/_102_ ),
    .B1(\lastadder/ksa32/_111_ ),
    .Y(\lastadder/ksa32/_112_ ));
 sky130_fd_sc_hd__xnor2_1 \lastadder/ksa32/_299_  (.A(\lastadder/ksa32/_110_ ),
    .B(\lastadder/ksa32/_112_ ),
    .Y(c[22]));
 sky130_fd_sc_hd__nor2_1 \lastadder/ksa32/_300_  (.A(_063_),
    .B(nextinp[23]),
    .Y(\lastadder/ksa32/_113_ ));
 sky130_fd_sc_hd__xor2_1 \lastadder/ksa32/_301_  (.A(_063_),
    .B(nextinp[23]),
    .X(\lastadder/ksa32/_114_ ));
 sky130_fd_sc_hd__nand2_1 \lastadder/ksa32/_302_  (.A(\lastadder/ksa32/_101_ ),
    .B(\lastadder/ksa32/_109_ ),
    .Y(\lastadder/ksa32/_115_ ));
 sky130_fd_sc_hd__o21ai_0 \lastadder/ksa32/_303_  (.A1(\lastadder/ksa32/_107_ ),
    .A2(\lastadder/ksa32/_115_ ),
    .B1(\lastadder/ksa32/_108_ ),
    .Y(\lastadder/ksa32/_116_ ));
 sky130_fd_sc_hd__o211a_1 \lastadder/ksa32/_304_  (.A1(\lastadder/ksa32/_107_ ),
    .A2(\lastadder/ksa32/_115_ ),
    .B1(\lastadder/ksa32/_114_ ),
    .C1(\lastadder/ksa32/_108_ ),
    .X(\lastadder/ksa32/_117_ ));
 sky130_fd_sc_hd__xnor2_1 \lastadder/ksa32/_305_  (.A(\lastadder/ksa32/_114_ ),
    .B(\lastadder/ksa32/_116_ ),
    .Y(c[23]));
 sky130_fd_sc_hd__xor2_1 \lastadder/ksa32/_306_  (.A(_064_),
    .B(nextinp[24]),
    .X(\lastadder/ksa32/_118_ ));
 sky130_fd_sc_hd__nand2_1 \lastadder/ksa32/_307_  (.A(\lastadder/ksa32/_110_ ),
    .B(\lastadder/ksa32/_114_ ),
    .Y(\lastadder/ksa32/_119_ ));
 sky130_fd_sc_hd__nor2_1 \lastadder/ksa32/_308_  (.A(\lastadder/ksa32/_109_ ),
    .B(\lastadder/ksa32/_113_ ),
    .Y(\lastadder/ksa32/_120_ ));
 sky130_fd_sc_hd__a21oi_1 \lastadder/ksa32/_309_  (.A1(_063_),
    .A2(nextinp[23]),
    .B1(\lastadder/ksa32/_120_ ),
    .Y(\lastadder/ksa32/_121_ ));
 sky130_fd_sc_hd__o21a_1 \lastadder/ksa32/_310_  (.A1(\lastadder/ksa32/_112_ ),
    .A2(\lastadder/ksa32/_119_ ),
    .B1(\lastadder/ksa32/_121_ ),
    .X(\lastadder/ksa32/_122_ ));
 sky130_fd_sc_hd__xnor2_1 \lastadder/ksa32/_311_  (.A(\lastadder/ksa32/_118_ ),
    .B(\lastadder/ksa32/_122_ ),
    .Y(c[24]));
 sky130_fd_sc_hd__nand2_1 \lastadder/ksa32/_312_  (.A(_065_),
    .B(nextinp[25]),
    .Y(\lastadder/ksa32/_123_ ));
 sky130_fd_sc_hd__xor2_1 \lastadder/ksa32/_313_  (.A(_065_),
    .B(nextinp[25]),
    .X(\lastadder/ksa32/_124_ ));
 sky130_fd_sc_hd__a22o_1 \lastadder/ksa32/_314_  (.A1(_063_),
    .A2(nextinp[23]),
    .B1(_064_),
    .B2(nextinp[24]),
    .X(\lastadder/ksa32/_125_ ));
 sky130_fd_sc_hd__o22ai_1 \lastadder/ksa32/_315_  (.A1(_064_),
    .A2(nextinp[24]),
    .B1(\lastadder/ksa32/_117_ ),
    .B2(\lastadder/ksa32/_125_ ),
    .Y(\lastadder/ksa32/_126_ ));
 sky130_fd_sc_hd__o221ai_1 \lastadder/ksa32/_316_  (.A1(_064_),
    .A2(nextinp[24]),
    .B1(\lastadder/ksa32/_117_ ),
    .B2(\lastadder/ksa32/_125_ ),
    .C1(\lastadder/ksa32/_124_ ),
    .Y(\lastadder/ksa32/_127_ ));
 sky130_fd_sc_hd__xnor2_1 \lastadder/ksa32/_317_  (.A(\lastadder/ksa32/_124_ ),
    .B(\lastadder/ksa32/_126_ ),
    .Y(c[25]));
 sky130_fd_sc_hd__o211ai_1 \lastadder/ksa32/_318_  (.A1(_065_),
    .A2(nextinp[25]),
    .B1(_064_),
    .C1(nextinp[24]),
    .Y(\lastadder/ksa32/_128_ ));
 sky130_fd_sc_hd__nand2_1 \lastadder/ksa32/_319_  (.A(\lastadder/ksa32/_118_ ),
    .B(\lastadder/ksa32/_124_ ),
    .Y(\lastadder/ksa32/_129_ ));
 sky130_fd_sc_hd__o211a_1 \lastadder/ksa32/_320_  (.A1(\lastadder/ksa32/_122_ ),
    .A2(\lastadder/ksa32/_129_ ),
    .B1(\lastadder/ksa32/_128_ ),
    .C1(\lastadder/ksa32/_123_ ),
    .X(\lastadder/ksa32/_130_ ));
 sky130_fd_sc_hd__nor2_1 \lastadder/ksa32/_321_  (.A(_066_),
    .B(nextinp[26]),
    .Y(\lastadder/ksa32/_131_ ));
 sky130_fd_sc_hd__nand2_1 \lastadder/ksa32/_322_  (.A(_066_),
    .B(nextinp[26]),
    .Y(\lastadder/ksa32/_132_ ));
 sky130_fd_sc_hd__nor2b_1 \lastadder/ksa32/_323_  (.A(\lastadder/ksa32/_131_ ),
    .B_N(\lastadder/ksa32/_132_ ),
    .Y(\lastadder/ksa32/_133_ ));
 sky130_fd_sc_hd__xnor2_1 \lastadder/ksa32/_324_  (.A(\lastadder/ksa32/_130_ ),
    .B(\lastadder/ksa32/_133_ ),
    .Y(c[26]));
 sky130_fd_sc_hd__nand2_1 \lastadder/ksa32/_325_  (.A(_067_),
    .B(nextinp[27]),
    .Y(\lastadder/ksa32/_134_ ));
 sky130_fd_sc_hd__xor2_1 \lastadder/ksa32/_326_  (.A(_067_),
    .B(nextinp[27]),
    .X(\lastadder/ksa32/_135_ ));
 sky130_fd_sc_hd__clkinv_1 \lastadder/ksa32/_327_  (.A(\lastadder/ksa32/_135_ ),
    .Y(\lastadder/ksa32/_136_ ));
 sky130_fd_sc_hd__a31oi_1 \lastadder/ksa32/_328_  (.A1(\lastadder/ksa32/_123_ ),
    .A2(\lastadder/ksa32/_127_ ),
    .A3(\lastadder/ksa32/_132_ ),
    .B1(\lastadder/ksa32/_131_ ),
    .Y(\lastadder/ksa32/_137_ ));
 sky130_fd_sc_hd__nor2_1 \lastadder/ksa32/_329_  (.A(\lastadder/ksa32/_135_ ),
    .B(\lastadder/ksa32/_137_ ),
    .Y(\lastadder/ksa32/_138_ ));
 sky130_fd_sc_hd__a311oi_1 \lastadder/ksa32/_330_  (.A1(\lastadder/ksa32/_123_ ),
    .A2(\lastadder/ksa32/_127_ ),
    .A3(\lastadder/ksa32/_132_ ),
    .B1(\lastadder/ksa32/_136_ ),
    .C1(\lastadder/ksa32/_131_ ),
    .Y(\lastadder/ksa32/_139_ ));
 sky130_fd_sc_hd__nor2_1 \lastadder/ksa32/_331_  (.A(\lastadder/ksa32/_138_ ),
    .B(\lastadder/ksa32/_139_ ),
    .Y(c[27]));
 sky130_fd_sc_hd__lpflow_inputiso1p_1 \lastadder/ksa32/_332_  (.A(_068_),
    .SLEEP(nextinp[28]),
    .X(\lastadder/ksa32/_140_ ));
 sky130_fd_sc_hd__nand2_1 \lastadder/ksa32/_333_  (.A(_068_),
    .B(nextinp[28]),
    .Y(\lastadder/ksa32/_141_ ));
 sky130_fd_sc_hd__nand2_1 \lastadder/ksa32/_334_  (.A(\lastadder/ksa32/_140_ ),
    .B(\lastadder/ksa32/_141_ ),
    .Y(\lastadder/ksa32/_142_ ));
 sky130_fd_sc_hd__nand2_1 \lastadder/ksa32/_335_  (.A(\lastadder/ksa32/_132_ ),
    .B(\lastadder/ksa32/_134_ ),
    .Y(\lastadder/ksa32/_143_ ));
 sky130_fd_sc_hd__o21ai_0 \lastadder/ksa32/_336_  (.A1(_067_),
    .A2(nextinp[27]),
    .B1(\lastadder/ksa32/_143_ ),
    .Y(\lastadder/ksa32/_144_ ));
 sky130_fd_sc_hd__nand2_1 \lastadder/ksa32/_337_  (.A(\lastadder/ksa32/_133_ ),
    .B(\lastadder/ksa32/_135_ ),
    .Y(\lastadder/ksa32/_145_ ));
 sky130_fd_sc_hd__o21ai_0 \lastadder/ksa32/_338_  (.A1(\lastadder/ksa32/_130_ ),
    .A2(\lastadder/ksa32/_145_ ),
    .B1(\lastadder/ksa32/_144_ ),
    .Y(\lastadder/ksa32/_146_ ));
 sky130_fd_sc_hd__xnor2_1 \lastadder/ksa32/_339_  (.A(\lastadder/ksa32/_142_ ),
    .B(\lastadder/ksa32/_146_ ),
    .Y(c[28]));
 sky130_fd_sc_hd__nor2_1 \lastadder/ksa32/_340_  (.A(_069_),
    .B(nextinp[29]),
    .Y(\lastadder/ksa32/_147_ ));
 sky130_fd_sc_hd__nand2_1 \lastadder/ksa32/_341_  (.A(_069_),
    .B(nextinp[29]),
    .Y(\lastadder/ksa32/_148_ ));
 sky130_fd_sc_hd__nor2b_1 \lastadder/ksa32/_342_  (.A(\lastadder/ksa32/_147_ ),
    .B_N(\lastadder/ksa32/_148_ ),
    .Y(\lastadder/ksa32/_149_ ));
 sky130_fd_sc_hd__nand2_1 \lastadder/ksa32/_343_  (.A(\lastadder/ksa32/_134_ ),
    .B(\lastadder/ksa32/_141_ ),
    .Y(\lastadder/ksa32/_150_ ));
 sky130_fd_sc_hd__o21ai_0 \lastadder/ksa32/_344_  (.A1(\lastadder/ksa32/_139_ ),
    .A2(\lastadder/ksa32/_150_ ),
    .B1(\lastadder/ksa32/_140_ ),
    .Y(\lastadder/ksa32/_151_ ));
 sky130_fd_sc_hd__o211ai_1 \lastadder/ksa32/_345_  (.A1(\lastadder/ksa32/_139_ ),
    .A2(\lastadder/ksa32/_150_ ),
    .B1(\lastadder/ksa32/_149_ ),
    .C1(\lastadder/ksa32/_140_ ),
    .Y(\lastadder/ksa32/_152_ ));
 sky130_fd_sc_hd__xnor2_1 \lastadder/ksa32/_346_  (.A(\lastadder/ksa32/_149_ ),
    .B(\lastadder/ksa32/_151_ ),
    .Y(c[29]));
 sky130_fd_sc_hd__o21ai_0 \lastadder/ksa32/_347_  (.A1(\lastadder/ksa32/_141_ ),
    .A2(\lastadder/ksa32/_147_ ),
    .B1(\lastadder/ksa32/_148_ ),
    .Y(\lastadder/ksa32/_153_ ));
 sky130_fd_sc_hd__a41oi_1 \lastadder/ksa32/_348_  (.A1(\lastadder/ksa32/_140_ ),
    .A2(\lastadder/ksa32/_141_ ),
    .A3(\lastadder/ksa32/_146_ ),
    .A4(\lastadder/ksa32/_149_ ),
    .B1(\lastadder/ksa32/_153_ ),
    .Y(\lastadder/ksa32/_154_ ));
 sky130_fd_sc_hd__nor2_1 \lastadder/ksa32/_349_  (.A(_070_),
    .B(nextinp[30]),
    .Y(\lastadder/ksa32/_155_ ));
 sky130_fd_sc_hd__nand2_1 \lastadder/ksa32/_350_  (.A(_070_),
    .B(nextinp[30]),
    .Y(\lastadder/ksa32/_156_ ));
 sky130_fd_sc_hd__nor2b_1 \lastadder/ksa32/_351_  (.A(\lastadder/ksa32/_155_ ),
    .B_N(\lastadder/ksa32/_156_ ),
    .Y(\lastadder/ksa32/_157_ ));
 sky130_fd_sc_hd__xnor2_1 \lastadder/ksa32/_352_  (.A(\lastadder/ksa32/_154_ ),
    .B(\lastadder/ksa32/_157_ ),
    .Y(c[30]));
 sky130_fd_sc_hd__nand2_1 \lastadder/ksa32/_353_  (.A(_071_),
    .B(nextinp[31]),
    .Y(\lastadder/ksa32/_158_ ));
 sky130_fd_sc_hd__xnor2_1 \lastadder/ksa32/_354_  (.A(_071_),
    .B(nextinp[31]),
    .Y(\lastadder/ksa32/_159_ ));
 sky130_fd_sc_hd__a31oi_1 \lastadder/ksa32/_355_  (.A1(\lastadder/ksa32/_148_ ),
    .A2(\lastadder/ksa32/_152_ ),
    .A3(\lastadder/ksa32/_156_ ),
    .B1(\lastadder/ksa32/_155_ ),
    .Y(\lastadder/ksa32/_160_ ));
 sky130_fd_sc_hd__xnor2_1 \lastadder/ksa32/_356_  (.A(\lastadder/ksa32/_159_ ),
    .B(\lastadder/ksa32/_160_ ),
    .Y(c[31]));
 sky130_fd_sc_hd__o211ai_1 \lastadder/ksa32/_357_  (.A1(\lastadder/ksa32/_154_ ),
    .A2(\lastadder/ksa32/_155_ ),
    .B1(\lastadder/ksa32/_156_ ),
    .C1(\lastadder/ksa32/_158_ ),
    .Y(\lastadder/ksa32/_161_ ));
 sky130_fd_sc_hd__o21a_1 \lastadder/ksa32/_358_  (.A1(_071_),
    .A2(nextinp[31]),
    .B1(\lastadder/ksa32/_161_ ),
    .X(\lastadder/Cout ));
 sky130_fd_sc_hd__conb_1 \v0/_35_  (.LO(\v0/_00_ ));
 sky130_fd_sc_hd__conb_1 \v0/_36_  (.LO(\v0/_01_ ));
 sky130_fd_sc_hd__conb_1 \v0/_37_  (.LO(\v0/_02_ ));
 sky130_fd_sc_hd__conb_1 \v0/_38_  (.LO(\v0/_03_ ));
 sky130_fd_sc_hd__conb_1 \v0/_39_  (.LO(\v0/_04_ ));
 sky130_fd_sc_hd__conb_1 \v0/_40_  (.LO(\v0/_05_ ));
 sky130_fd_sc_hd__conb_1 \v0/_41_  (.LO(\v0/_06_ ));
 sky130_fd_sc_hd__conb_1 \v0/_42_  (.LO(\v0/_07_ ));
 sky130_fd_sc_hd__conb_1 \v0/_43_  (.LO(\v0/_08_ ));
 sky130_fd_sc_hd__conb_1 \v0/_44_  (.LO(\v0/_09_ ));
 sky130_fd_sc_hd__conb_1 \v0/_45_  (.LO(\v0/_10_ ));
 sky130_fd_sc_hd__conb_1 \v0/_46_  (.LO(\v0/_11_ ));
 sky130_fd_sc_hd__conb_1 \v0/_47_  (.LO(\v0/_12_ ));
 sky130_fd_sc_hd__conb_1 \v0/_48_  (.LO(\v0/_13_ ));
 sky130_fd_sc_hd__conb_1 \v0/_49_  (.LO(\v0/_14_ ));
 sky130_fd_sc_hd__conb_1 \v0/_50_  (.LO(\v0/_15_ ));
 sky130_fd_sc_hd__conb_1 \v0/_51_  (.LO(\v0/_16_ ));
 sky130_fd_sc_hd__conb_1 \v0/_52_  (.LO(\v0/_17_ ));
 sky130_fd_sc_hd__conb_1 \v0/_53_  (.LO(\v0/_18_ ));
 sky130_fd_sc_hd__conb_1 \v0/_54_  (.LO(\v0/_19_ ));
 sky130_fd_sc_hd__conb_1 \v0/_55_  (.LO(\v0/_20_ ));
 sky130_fd_sc_hd__conb_1 \v0/_56_  (.LO(\v0/_21_ ));
 sky130_fd_sc_hd__conb_1 \v0/_57_  (.LO(\v0/_22_ ));
 sky130_fd_sc_hd__conb_1 \v0/_58_  (.LO(\v0/_23_ ));
 sky130_fd_sc_hd__conb_1 \v0/_59_  (.LO(\v0/_24_ ));
 sky130_fd_sc_hd__conb_1 \v0/_60_  (.LO(\v0/_25_ ));
 sky130_fd_sc_hd__conb_1 \v0/_61_  (.LO(\v0/_26_ ));
 sky130_fd_sc_hd__conb_1 \v0/_62_  (.LO(\v0/_27_ ));
 sky130_fd_sc_hd__conb_1 \v0/_63_  (.LO(\v0/_28_ ));
 sky130_fd_sc_hd__conb_1 \v0/_64_  (.LO(\v0/_29_ ));
 sky130_fd_sc_hd__conb_1 \v0/_65_  (.LO(\v0/_30_ ));
 sky130_fd_sc_hd__conb_1 \v0/_66_  (.LO(\v0/_31_ ));
 sky130_fd_sc_hd__conb_1 \v0/_67_  (.LO(\v0/_32_ ));
 sky130_fd_sc_hd__conb_1 \v0/_68_  (.LO(\v0/_33_ ));
 sky130_fd_sc_hd__conb_1 \v0/_69_  (.LO(\v0/_34_ ));
 sky130_fd_sc_hd__conb_1 \v0/z1/_19_  (.LO(\v0/z1/_00_ ));
 sky130_fd_sc_hd__conb_1 \v0/z1/_20_  (.LO(\v0/z1/_01_ ));
 sky130_fd_sc_hd__conb_1 \v0/z1/_21_  (.LO(\v0/z1/_02_ ));
 sky130_fd_sc_hd__conb_1 \v0/z1/_22_  (.LO(\v0/z1/_03_ ));
 sky130_fd_sc_hd__conb_1 \v0/z1/_23_  (.LO(\v0/z1/_04_ ));
 sky130_fd_sc_hd__conb_1 \v0/z1/_24_  (.LO(\v0/z1/_05_ ));
 sky130_fd_sc_hd__conb_1 \v0/z1/_25_  (.LO(\v0/z1/_06_ ));
 sky130_fd_sc_hd__conb_1 \v0/z1/_26_  (.LO(\v0/z1/_07_ ));
 sky130_fd_sc_hd__conb_1 \v0/z1/_27_  (.LO(\v0/z1/_08_ ));
 sky130_fd_sc_hd__conb_1 \v0/z1/_28_  (.LO(\v0/z1/_09_ ));
 sky130_fd_sc_hd__conb_1 \v0/z1/_29_  (.LO(\v0/z1/_10_ ));
 sky130_fd_sc_hd__conb_1 \v0/z1/_30_  (.LO(\v0/z1/_11_ ));
 sky130_fd_sc_hd__conb_1 \v0/z1/_31_  (.LO(\v0/z1/_12_ ));
 sky130_fd_sc_hd__conb_1 \v0/z1/_32_  (.LO(\v0/z1/_13_ ));
 sky130_fd_sc_hd__conb_1 \v0/z1/_33_  (.LO(\v0/z1/_14_ ));
 sky130_fd_sc_hd__conb_1 \v0/z1/_34_  (.LO(\v0/z1/_15_ ));
 sky130_fd_sc_hd__conb_1 \v0/z1/_35_  (.LO(\v0/z1/_16_ ));
 sky130_fd_sc_hd__conb_1 \v0/z1/_36_  (.LO(\v0/z1/_17_ ));
 sky130_fd_sc_hd__conb_1 \v0/z1/_37_  (.LO(\v0/z1/_18_ ));
 sky130_fd_sc_hd__conb_1 \v0/z1/z1/_11_  (.LO(\v0/z1/z1/_00_ ));
 sky130_fd_sc_hd__conb_1 \v0/z1/z1/_12_  (.LO(\v0/z1/z1/_01_ ));
 sky130_fd_sc_hd__conb_1 \v0/z1/z1/_13_  (.LO(\v0/z1/z1/_02_ ));
 sky130_fd_sc_hd__conb_1 \v0/z1/z1/_14_  (.LO(\v0/z1/z1/_03_ ));
 sky130_fd_sc_hd__conb_1 \v0/z1/z1/_15_  (.LO(\v0/z1/z1/_04_ ));
 sky130_fd_sc_hd__conb_1 \v0/z1/z1/_16_  (.LO(\v0/z1/z1/_05_ ));
 sky130_fd_sc_hd__conb_1 \v0/z1/z1/_17_  (.LO(\v0/z1/z1/_06_ ));
 sky130_fd_sc_hd__conb_1 \v0/z1/z1/_18_  (.LO(\v0/z1/z1/_07_ ));
 sky130_fd_sc_hd__conb_1 \v0/z1/z1/_19_  (.LO(\v0/z1/z1/_08_ ));
 sky130_fd_sc_hd__conb_1 \v0/z1/z1/_20_  (.LO(\v0/z1/z1/_09_ ));
 sky130_fd_sc_hd__conb_1 \v0/z1/z1/_21_  (.LO(\v0/z1/z1/_10_ ));
 sky130_fd_sc_hd__and2_0 \v0/z1/z1/z1/_0_  (.A(b[0]),
    .B(a[0]),
    .X(unsign[0]));
 sky130_fd_sc_hd__and2_0 \v0/z1/z1/z1/_1_  (.A(b[0]),
    .B(abs_a[1]),
    .X(\v0/z1/z1/z1/temp [0]));
 sky130_fd_sc_hd__and2_0 \v0/z1/z1/z1/_2_  (.A(a[0]),
    .B(abs_b[1]),
    .X(\v0/z1/z1/z1/temp [1]));
 sky130_fd_sc_hd__and2_0 \v0/z1/z1/z1/_3_  (.A(abs_a[1]),
    .B(abs_b[1]),
    .X(\v0/z1/z1/z1/temp [2]));
 sky130_fd_sc_hd__and2_0 \v0/z1/z1/z1/z1/_0_  (.A(\v0/z1/z1/z1/temp [1]),
    .B(\v0/z1/z1/z1/temp [0]),
    .X(\v0/z1/z1/z1/temp [3]));
 sky130_fd_sc_hd__xor2_1 \v0/z1/z1/z1/z1/_1_  (.A(\v0/z1/z1/z1/temp [1]),
    .B(\v0/z1/z1/z1/temp [0]),
    .X(unsign[1]));
 sky130_fd_sc_hd__and2_0 \v0/z1/z1/z1/z2/_0_  (.A(\v0/z1/z1/z1/temp [3]),
    .B(\v0/z1/z1/z1/temp [2]),
    .X(\v0/z1/z1/q0 [3]));
 sky130_fd_sc_hd__xor2_1 \v0/z1/z1/z1/z2/_1_  (.A(\v0/z1/z1/z1/temp [3]),
    .B(\v0/z1/z1/z1/temp [2]),
    .X(\v0/z1/z1/q0 [2]));
 sky130_fd_sc_hd__and2_0 \v0/z1/z1/z2/_0_  (.A(b[0]),
    .B(abs_a[2]),
    .X(\v0/z1/z1/q1 [0]));
 sky130_fd_sc_hd__and2_0 \v0/z1/z1/z2/_1_  (.A(b[0]),
    .B(abs_a[3]),
    .X(\v0/z1/z1/z2/temp [0]));
 sky130_fd_sc_hd__and2_0 \v0/z1/z1/z2/_2_  (.A(abs_a[2]),
    .B(abs_b[1]),
    .X(\v0/z1/z1/z2/temp [1]));
 sky130_fd_sc_hd__and2_0 \v0/z1/z1/z2/_3_  (.A(abs_a[3]),
    .B(abs_b[1]),
    .X(\v0/z1/z1/z2/temp [2]));
 sky130_fd_sc_hd__and2_0 \v0/z1/z1/z2/z1/_0_  (.A(\v0/z1/z1/z2/temp [1]),
    .B(\v0/z1/z1/z2/temp [0]),
    .X(\v0/z1/z1/z2/temp [3]));
 sky130_fd_sc_hd__xor2_1 \v0/z1/z1/z2/z1/_1_  (.A(\v0/z1/z1/z2/temp [1]),
    .B(\v0/z1/z1/z2/temp [0]),
    .X(\v0/z1/z1/q1 [1]));
 sky130_fd_sc_hd__and2_0 \v0/z1/z1/z2/z2/_0_  (.A(\v0/z1/z1/z2/temp [3]),
    .B(\v0/z1/z1/z2/temp [2]),
    .X(\v0/z1/z1/q1 [3]));
 sky130_fd_sc_hd__xor2_1 \v0/z1/z1/z2/z2/_1_  (.A(\v0/z1/z1/z2/temp [3]),
    .B(\v0/z1/z1/z2/temp [2]),
    .X(\v0/z1/z1/q1 [2]));
 sky130_fd_sc_hd__and2_0 \v0/z1/z1/z3/_0_  (.A(abs_b[2]),
    .B(a[0]),
    .X(\v0/z1/z1/q2 [0]));
 sky130_fd_sc_hd__and2_0 \v0/z1/z1/z3/_1_  (.A(abs_b[2]),
    .B(abs_a[1]),
    .X(\v0/z1/z1/z3/temp [0]));
 sky130_fd_sc_hd__and2_0 \v0/z1/z1/z3/_2_  (.A(a[0]),
    .B(abs_b[3]),
    .X(\v0/z1/z1/z3/temp [1]));
 sky130_fd_sc_hd__and2_0 \v0/z1/z1/z3/_3_  (.A(abs_a[1]),
    .B(abs_b[3]),
    .X(\v0/z1/z1/z3/temp [2]));
 sky130_fd_sc_hd__and2_0 \v0/z1/z1/z3/z1/_0_  (.A(\v0/z1/z1/z3/temp [1]),
    .B(\v0/z1/z1/z3/temp [0]),
    .X(\v0/z1/z1/z3/temp [3]));
 sky130_fd_sc_hd__xor2_1 \v0/z1/z1/z3/z1/_1_  (.A(\v0/z1/z1/z3/temp [1]),
    .B(\v0/z1/z1/z3/temp [0]),
    .X(\v0/z1/z1/q2 [1]));
 sky130_fd_sc_hd__and2_0 \v0/z1/z1/z3/z2/_0_  (.A(\v0/z1/z1/z3/temp [3]),
    .B(\v0/z1/z1/z3/temp [2]),
    .X(\v0/z1/z1/q2 [3]));
 sky130_fd_sc_hd__xor2_1 \v0/z1/z1/z3/z2/_1_  (.A(\v0/z1/z1/z3/temp [3]),
    .B(\v0/z1/z1/z3/temp [2]),
    .X(\v0/z1/z1/q2 [2]));
 sky130_fd_sc_hd__and2_0 \v0/z1/z1/z4/_0_  (.A(abs_b[2]),
    .B(abs_a[2]),
    .X(\v0/z1/z1/q3 [0]));
 sky130_fd_sc_hd__and2_0 \v0/z1/z1/z4/_1_  (.A(abs_b[2]),
    .B(abs_a[3]),
    .X(\v0/z1/z1/z4/temp [0]));
 sky130_fd_sc_hd__and2_0 \v0/z1/z1/z4/_2_  (.A(abs_a[2]),
    .B(abs_b[3]),
    .X(\v0/z1/z1/z4/temp [1]));
 sky130_fd_sc_hd__and2_0 \v0/z1/z1/z4/_3_  (.A(abs_a[3]),
    .B(abs_b[3]),
    .X(\v0/z1/z1/z4/temp [2]));
 sky130_fd_sc_hd__and2_0 \v0/z1/z1/z4/z1/_0_  (.A(\v0/z1/z1/z4/temp [1]),
    .B(\v0/z1/z1/z4/temp [0]),
    .X(\v0/z1/z1/z4/temp [3]));
 sky130_fd_sc_hd__xor2_1 \v0/z1/z1/z4/z1/_1_  (.A(\v0/z1/z1/z4/temp [1]),
    .B(\v0/z1/z1/z4/temp [0]),
    .X(\v0/z1/z1/q3 [1]));
 sky130_fd_sc_hd__and2_0 \v0/z1/z1/z4/z2/_0_  (.A(\v0/z1/z1/z4/temp [3]),
    .B(\v0/z1/z1/z4/temp [2]),
    .X(\v0/z1/z1/q3 [3]));
 sky130_fd_sc_hd__xor2_1 \v0/z1/z1/z4/z2/_1_  (.A(\v0/z1/z1/z4/temp [3]),
    .B(\v0/z1/z1/z4/temp [2]),
    .X(\v0/z1/z1/q3 [2]));
 sky130_fd_sc_hd__xnor2_1 \v0/z1/z1/z5/_07_  (.A(\v0/z1/z1/q0 [2]),
    .B(\v0/z1/z1/q1 [0]),
    .Y(\v0/z1/z1/z5/_00_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z1/z1/z5/_08_  (.A(\v0/z1/z1/_02_ ),
    .B(\v0/z1/z1/z5/_00_ ),
    .Y(\v0/z1/z1/q4 [0]));
 sky130_fd_sc_hd__maj3_1 \v0/z1/z1/z5/_09_  (.A(\v0/z1/z1/q0 [2]),
    .B(\v0/z1/z1/q1 [0]),
    .C(\v0/z1/z1/_02_ ),
    .X(\v0/z1/z1/z5/_01_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z1/z1/z5/_10_  (.A(\v0/z1/z1/q0 [3]),
    .B(\v0/z1/z1/q1 [1]),
    .Y(\v0/z1/z1/z5/_02_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z1/z1/z5/_11_  (.A(\v0/z1/z1/z5/_01_ ),
    .B(\v0/z1/z1/z5/_02_ ),
    .Y(\v0/z1/z1/q4 [1]));
 sky130_fd_sc_hd__maj3_1 \v0/z1/z1/z5/_12_  (.A(\v0/z1/z1/q0 [3]),
    .B(\v0/z1/z1/q1 [1]),
    .C(\v0/z1/z1/z5/_01_ ),
    .X(\v0/z1/z1/z5/_03_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z1/z1/z5/_13_  (.A(\v0/z1/z1/_00_ ),
    .B(\v0/z1/z1/q1 [2]),
    .Y(\v0/z1/z1/z5/_04_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z1/z1/z5/_14_  (.A(\v0/z1/z1/z5/_03_ ),
    .B(\v0/z1/z1/z5/_04_ ),
    .Y(\v0/z1/z1/q4 [2]));
 sky130_fd_sc_hd__maj3_1 \v0/z1/z1/z5/_15_  (.A(\v0/z1/z1/_00_ ),
    .B(\v0/z1/z1/q1 [2]),
    .C(\v0/z1/z1/z5/_03_ ),
    .X(\v0/z1/z1/z5/_05_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z1/z1/z5/_16_  (.A(\v0/z1/z1/_01_ ),
    .B(\v0/z1/z1/q1 [3]),
    .Y(\v0/z1/z1/z5/_06_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z1/z1/z5/_17_  (.A(\v0/z1/z1/z5/_05_ ),
    .B(\v0/z1/z1/z5/_06_ ),
    .Y(\v0/z1/z1/q4 [3]));
 sky130_fd_sc_hd__maj3_1 \v0/z1/z1/z5/_18_  (.A(\v0/z1/z1/_01_ ),
    .B(\v0/z1/z1/q1 [3]),
    .C(\v0/z1/z1/z5/_05_ ),
    .X(\v0/z1/z1/z5/Cout ));
 sky130_fd_sc_hd__xnor2_1 \v0/z1/z1/z6/_19_  (.A(\v0/z1/z1/_05_ ),
    .B(\v0/z1/z1/q2 [0]),
    .Y(\v0/z1/z1/z6/_00_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z1/z1/z6/_20_  (.A(\v0/z1/z1/_07_ ),
    .B(\v0/z1/z1/z6/_00_ ),
    .Y(\v0/z1/z1/q5 [0]));
 sky130_fd_sc_hd__maj3_1 \v0/z1/z1/z6/_21_  (.A(\v0/z1/z1/_05_ ),
    .B(\v0/z1/z1/q2 [0]),
    .C(\v0/z1/z1/_07_ ),
    .X(\v0/z1/z1/z6/_01_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z1/z1/z6/_22_  (.A(\v0/z1/z1/_06_ ),
    .B(\v0/z1/z1/q2 [1]),
    .Y(\v0/z1/z1/z6/_02_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z1/z1/z6/_23_  (.A(\v0/z1/z1/z6/_01_ ),
    .B(\v0/z1/z1/z6/_02_ ),
    .Y(\v0/z1/z1/q5 [1]));
 sky130_fd_sc_hd__maj3_1 \v0/z1/z1/z6/_24_  (.A(\v0/z1/z1/_06_ ),
    .B(\v0/z1/z1/q2 [1]),
    .C(\v0/z1/z1/z6/_01_ ),
    .X(\v0/z1/z1/z6/_03_ ));
 sky130_fd_sc_hd__lpflow_inputiso1p_1 \v0/z1/z1/z6/_25_  (.A(\v0/z1/z1/q3 [0]),
    .SLEEP(\v0/z1/z1/q2 [2]),
    .X(\v0/z1/z1/z6/_04_ ));
 sky130_fd_sc_hd__and2_0 \v0/z1/z1/z6/_26_  (.A(\v0/z1/z1/q3 [0]),
    .B(\v0/z1/z1/q2 [2]),
    .X(\v0/z1/z1/z6/_05_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z1/z1/z6/_27_  (.A(\v0/z1/z1/q3 [0]),
    .B(\v0/z1/z1/q2 [2]),
    .Y(\v0/z1/z1/z6/_06_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z1/z1/z6/_28_  (.A(\v0/z1/z1/z6/_04_ ),
    .B(\v0/z1/z1/z6/_06_ ),
    .Y(\v0/z1/z1/z6/_07_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z1/z1/z6/_29_  (.A(\v0/z1/z1/z6/_03_ ),
    .B(\v0/z1/z1/z6/_07_ ),
    .Y(\v0/z1/z1/q5 [2]));
 sky130_fd_sc_hd__nand2_1 \v0/z1/z1/z6/_30_  (.A(\v0/z1/z1/q3 [1]),
    .B(\v0/z1/z1/q2 [3]),
    .Y(\v0/z1/z1/z6/_08_ ));
 sky130_fd_sc_hd__xor2_1 \v0/z1/z1/z6/_31_  (.A(\v0/z1/z1/q3 [1]),
    .B(\v0/z1/z1/q2 [3]),
    .X(\v0/z1/z1/z6/_09_ ));
 sky130_fd_sc_hd__o21ai_0 \v0/z1/z1/z6/_32_  (.A1(\v0/z1/z1/z6/_03_ ),
    .A2(\v0/z1/z1/z6/_05_ ),
    .B1(\v0/z1/z1/z6/_04_ ),
    .Y(\v0/z1/z1/z6/_10_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z1/z1/z6/_33_  (.A(\v0/z1/z1/z6/_09_ ),
    .B(\v0/z1/z1/z6/_10_ ),
    .Y(\v0/z1/z1/q5 [3]));
 sky130_fd_sc_hd__nor2_1 \v0/z1/z1/z6/_34_  (.A(\v0/z1/z1/q3 [2]),
    .B(\v0/z1/z1/_03_ ),
    .Y(\v0/z1/z1/z6/_11_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z1/z1/z6/_35_  (.A(\v0/z1/z1/q3 [2]),
    .B(\v0/z1/z1/_03_ ),
    .Y(\v0/z1/z1/z6/_12_ ));
 sky130_fd_sc_hd__nand2b_1 \v0/z1/z1/z6/_36_  (.A_N(\v0/z1/z1/z6/_11_ ),
    .B(\v0/z1/z1/z6/_12_ ),
    .Y(\v0/z1/z1/z6/_13_ ));
 sky130_fd_sc_hd__o221ai_1 \v0/z1/z1/z6/_37_  (.A1(\v0/z1/z1/q3 [1]),
    .A2(\v0/z1/z1/q2 [3]),
    .B1(\v0/z1/z1/z6/_03_ ),
    .B2(\v0/z1/z1/z6/_05_ ),
    .C1(\v0/z1/z1/z6/_04_ ),
    .Y(\v0/z1/z1/z6/_14_ ));
 sky130_fd_sc_hd__a21oi_1 \v0/z1/z1/z6/_38_  (.A1(\v0/z1/z1/z6/_08_ ),
    .A2(\v0/z1/z1/z6/_14_ ),
    .B1(\v0/z1/z1/z6/_13_ ),
    .Y(\v0/z1/z1/z6/_15_ ));
 sky130_fd_sc_hd__and3_1 \v0/z1/z1/z6/_39_  (.A(\v0/z1/z1/z6/_08_ ),
    .B(\v0/z1/z1/z6/_13_ ),
    .C(\v0/z1/z1/z6/_14_ ),
    .X(\v0/z1/z1/z6/_16_ ));
 sky130_fd_sc_hd__nor2_1 \v0/z1/z1/z6/_40_  (.A(\v0/z1/z1/z6/_15_ ),
    .B(\v0/z1/z1/z6/_16_ ),
    .Y(\v0/z1/z1/q5 [4]));
 sky130_fd_sc_hd__xnor2_1 \v0/z1/z1/z6/_41_  (.A(\v0/z1/z1/q3 [3]),
    .B(\v0/z1/z1/_04_ ),
    .Y(\v0/z1/z1/z6/_17_ ));
 sky130_fd_sc_hd__a31oi_1 \v0/z1/z1/z6/_42_  (.A1(\v0/z1/z1/z6/_08_ ),
    .A2(\v0/z1/z1/z6/_12_ ),
    .A3(\v0/z1/z1/z6/_14_ ),
    .B1(\v0/z1/z1/z6/_11_ ),
    .Y(\v0/z1/z1/z6/_18_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z1/z1/z6/_43_  (.A(\v0/z1/z1/z6/_17_ ),
    .B(\v0/z1/z1/z6/_18_ ),
    .Y(\v0/z1/z1/q5 [5]));
 sky130_fd_sc_hd__maj3_1 \v0/z1/z1/z6/_44_  (.A(\v0/z1/z1/q3 [3]),
    .B(\v0/z1/z1/_04_ ),
    .C(\v0/z1/z1/z6/_18_ ),
    .X(\v0/z1/z1/z6/Cout ));
 sky130_fd_sc_hd__xnor2_1 \v0/z1/z1/z7/_19_  (.A(\v0/z1/z1/q5 [0]),
    .B(\v0/z1/z1/q4 [0]),
    .Y(\v0/z1/z1/z7/_00_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z1/z1/z7/_20_  (.A(\v0/z1/z1/_10_ ),
    .B(\v0/z1/z1/z7/_00_ ),
    .Y(unsign[2]));
 sky130_fd_sc_hd__maj3_1 \v0/z1/z1/z7/_21_  (.A(\v0/z1/z1/q5 [0]),
    .B(\v0/z1/z1/q4 [0]),
    .C(\v0/z1/z1/_10_ ),
    .X(\v0/z1/z1/z7/_01_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z1/z1/z7/_22_  (.A(\v0/z1/z1/q5 [1]),
    .B(\v0/z1/z1/q4 [1]),
    .Y(\v0/z1/z1/z7/_02_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z1/z1/z7/_23_  (.A(\v0/z1/z1/z7/_01_ ),
    .B(\v0/z1/z1/z7/_02_ ),
    .Y(unsign[3]));
 sky130_fd_sc_hd__maj3_1 \v0/z1/z1/z7/_24_  (.A(\v0/z1/z1/q5 [1]),
    .B(\v0/z1/z1/q4 [1]),
    .C(\v0/z1/z1/z7/_01_ ),
    .X(\v0/z1/z1/z7/_03_ ));
 sky130_fd_sc_hd__lpflow_inputiso1p_1 \v0/z1/z1/z7/_25_  (.A(\v0/z1/z1/q5 [2]),
    .SLEEP(\v0/z1/z1/q4 [2]),
    .X(\v0/z1/z1/z7/_04_ ));
 sky130_fd_sc_hd__and2_0 \v0/z1/z1/z7/_26_  (.A(\v0/z1/z1/q5 [2]),
    .B(\v0/z1/z1/q4 [2]),
    .X(\v0/z1/z1/z7/_05_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z1/z1/z7/_27_  (.A(\v0/z1/z1/q5 [2]),
    .B(\v0/z1/z1/q4 [2]),
    .Y(\v0/z1/z1/z7/_06_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z1/z1/z7/_28_  (.A(\v0/z1/z1/z7/_04_ ),
    .B(\v0/z1/z1/z7/_06_ ),
    .Y(\v0/z1/z1/z7/_07_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z1/z1/z7/_29_  (.A(\v0/z1/z1/z7/_03_ ),
    .B(\v0/z1/z1/z7/_07_ ),
    .Y(\v0/z1/q0 [4]));
 sky130_fd_sc_hd__nand2_1 \v0/z1/z1/z7/_30_  (.A(\v0/z1/z1/q5 [3]),
    .B(\v0/z1/z1/q4 [3]),
    .Y(\v0/z1/z1/z7/_08_ ));
 sky130_fd_sc_hd__xor2_1 \v0/z1/z1/z7/_31_  (.A(\v0/z1/z1/q5 [3]),
    .B(\v0/z1/z1/q4 [3]),
    .X(\v0/z1/z1/z7/_09_ ));
 sky130_fd_sc_hd__o21ai_0 \v0/z1/z1/z7/_32_  (.A1(\v0/z1/z1/z7/_03_ ),
    .A2(\v0/z1/z1/z7/_05_ ),
    .B1(\v0/z1/z1/z7/_04_ ),
    .Y(\v0/z1/z1/z7/_10_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z1/z1/z7/_33_  (.A(\v0/z1/z1/z7/_09_ ),
    .B(\v0/z1/z1/z7/_10_ ),
    .Y(\v0/z1/q0 [5]));
 sky130_fd_sc_hd__nor2_1 \v0/z1/z1/z7/_34_  (.A(\v0/z1/z1/q5 [4]),
    .B(\v0/z1/z1/_08_ ),
    .Y(\v0/z1/z1/z7/_11_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z1/z1/z7/_35_  (.A(\v0/z1/z1/q5 [4]),
    .B(\v0/z1/z1/_08_ ),
    .Y(\v0/z1/z1/z7/_12_ ));
 sky130_fd_sc_hd__nand2b_1 \v0/z1/z1/z7/_36_  (.A_N(\v0/z1/z1/z7/_11_ ),
    .B(\v0/z1/z1/z7/_12_ ),
    .Y(\v0/z1/z1/z7/_13_ ));
 sky130_fd_sc_hd__o221ai_1 \v0/z1/z1/z7/_37_  (.A1(\v0/z1/z1/q5 [3]),
    .A2(\v0/z1/z1/q4 [3]),
    .B1(\v0/z1/z1/z7/_03_ ),
    .B2(\v0/z1/z1/z7/_05_ ),
    .C1(\v0/z1/z1/z7/_04_ ),
    .Y(\v0/z1/z1/z7/_14_ ));
 sky130_fd_sc_hd__a21oi_1 \v0/z1/z1/z7/_38_  (.A1(\v0/z1/z1/z7/_08_ ),
    .A2(\v0/z1/z1/z7/_14_ ),
    .B1(\v0/z1/z1/z7/_13_ ),
    .Y(\v0/z1/z1/z7/_15_ ));
 sky130_fd_sc_hd__and3_1 \v0/z1/z1/z7/_39_  (.A(\v0/z1/z1/z7/_08_ ),
    .B(\v0/z1/z1/z7/_13_ ),
    .C(\v0/z1/z1/z7/_14_ ),
    .X(\v0/z1/z1/z7/_16_ ));
 sky130_fd_sc_hd__nor2_1 \v0/z1/z1/z7/_40_  (.A(\v0/z1/z1/z7/_15_ ),
    .B(\v0/z1/z1/z7/_16_ ),
    .Y(\v0/z1/q0 [6]));
 sky130_fd_sc_hd__xnor2_1 \v0/z1/z1/z7/_41_  (.A(\v0/z1/z1/q5 [5]),
    .B(\v0/z1/z1/_09_ ),
    .Y(\v0/z1/z1/z7/_17_ ));
 sky130_fd_sc_hd__a31oi_1 \v0/z1/z1/z7/_42_  (.A1(\v0/z1/z1/z7/_08_ ),
    .A2(\v0/z1/z1/z7/_12_ ),
    .A3(\v0/z1/z1/z7/_14_ ),
    .B1(\v0/z1/z1/z7/_11_ ),
    .Y(\v0/z1/z1/z7/_18_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z1/z1/z7/_43_  (.A(\v0/z1/z1/z7/_17_ ),
    .B(\v0/z1/z1/z7/_18_ ),
    .Y(\v0/z1/q0 [7]));
 sky130_fd_sc_hd__maj3_1 \v0/z1/z1/z7/_44_  (.A(\v0/z1/z1/q5 [5]),
    .B(\v0/z1/z1/_09_ ),
    .C(\v0/z1/z1/z7/_18_ ),
    .X(\v0/z1/z1/z7/Cout ));
 sky130_fd_sc_hd__conb_1 \v0/z1/z2/_11_  (.LO(\v0/z1/z2/_00_ ));
 sky130_fd_sc_hd__conb_1 \v0/z1/z2/_12_  (.LO(\v0/z1/z2/_01_ ));
 sky130_fd_sc_hd__conb_1 \v0/z1/z2/_13_  (.LO(\v0/z1/z2/_02_ ));
 sky130_fd_sc_hd__conb_1 \v0/z1/z2/_14_  (.LO(\v0/z1/z2/_03_ ));
 sky130_fd_sc_hd__conb_1 \v0/z1/z2/_15_  (.LO(\v0/z1/z2/_04_ ));
 sky130_fd_sc_hd__conb_1 \v0/z1/z2/_16_  (.LO(\v0/z1/z2/_05_ ));
 sky130_fd_sc_hd__conb_1 \v0/z1/z2/_17_  (.LO(\v0/z1/z2/_06_ ));
 sky130_fd_sc_hd__conb_1 \v0/z1/z2/_18_  (.LO(\v0/z1/z2/_07_ ));
 sky130_fd_sc_hd__conb_1 \v0/z1/z2/_19_  (.LO(\v0/z1/z2/_08_ ));
 sky130_fd_sc_hd__conb_1 \v0/z1/z2/_20_  (.LO(\v0/z1/z2/_09_ ));
 sky130_fd_sc_hd__conb_1 \v0/z1/z2/_21_  (.LO(\v0/z1/z2/_10_ ));
 sky130_fd_sc_hd__and2_0 \v0/z1/z2/z1/_0_  (.A(b[0]),
    .B(abs_a[4]),
    .X(\v0/z1/q1 [0]));
 sky130_fd_sc_hd__and2_0 \v0/z1/z2/z1/_1_  (.A(b[0]),
    .B(abs_a[5]),
    .X(\v0/z1/z2/z1/temp [0]));
 sky130_fd_sc_hd__and2_0 \v0/z1/z2/z1/_2_  (.A(abs_a[4]),
    .B(abs_b[1]),
    .X(\v0/z1/z2/z1/temp [1]));
 sky130_fd_sc_hd__and2_0 \v0/z1/z2/z1/_3_  (.A(abs_a[5]),
    .B(abs_b[1]),
    .X(\v0/z1/z2/z1/temp [2]));
 sky130_fd_sc_hd__and2_0 \v0/z1/z2/z1/z1/_0_  (.A(\v0/z1/z2/z1/temp [1]),
    .B(\v0/z1/z2/z1/temp [0]),
    .X(\v0/z1/z2/z1/temp [3]));
 sky130_fd_sc_hd__xor2_1 \v0/z1/z2/z1/z1/_1_  (.A(\v0/z1/z2/z1/temp [1]),
    .B(\v0/z1/z2/z1/temp [0]),
    .X(\v0/z1/q1 [1]));
 sky130_fd_sc_hd__and2_0 \v0/z1/z2/z1/z2/_0_  (.A(\v0/z1/z2/z1/temp [3]),
    .B(\v0/z1/z2/z1/temp [2]),
    .X(\v0/z1/z2/q0 [3]));
 sky130_fd_sc_hd__xor2_1 \v0/z1/z2/z1/z2/_1_  (.A(\v0/z1/z2/z1/temp [3]),
    .B(\v0/z1/z2/z1/temp [2]),
    .X(\v0/z1/z2/q0 [2]));
 sky130_fd_sc_hd__and2_0 \v0/z1/z2/z2/_0_  (.A(b[0]),
    .B(abs_a[6]),
    .X(\v0/z1/z2/q1 [0]));
 sky130_fd_sc_hd__and2_0 \v0/z1/z2/z2/_1_  (.A(b[0]),
    .B(abs_a[7]),
    .X(\v0/z1/z2/z2/temp [0]));
 sky130_fd_sc_hd__and2_0 \v0/z1/z2/z2/_2_  (.A(abs_a[6]),
    .B(abs_b[1]),
    .X(\v0/z1/z2/z2/temp [1]));
 sky130_fd_sc_hd__and2_0 \v0/z1/z2/z2/_3_  (.A(abs_a[7]),
    .B(abs_b[1]),
    .X(\v0/z1/z2/z2/temp [2]));
 sky130_fd_sc_hd__and2_0 \v0/z1/z2/z2/z1/_0_  (.A(\v0/z1/z2/z2/temp [1]),
    .B(\v0/z1/z2/z2/temp [0]),
    .X(\v0/z1/z2/z2/temp [3]));
 sky130_fd_sc_hd__xor2_1 \v0/z1/z2/z2/z1/_1_  (.A(\v0/z1/z2/z2/temp [1]),
    .B(\v0/z1/z2/z2/temp [0]),
    .X(\v0/z1/z2/q1 [1]));
 sky130_fd_sc_hd__and2_0 \v0/z1/z2/z2/z2/_0_  (.A(\v0/z1/z2/z2/temp [3]),
    .B(\v0/z1/z2/z2/temp [2]),
    .X(\v0/z1/z2/q1 [3]));
 sky130_fd_sc_hd__xor2_1 \v0/z1/z2/z2/z2/_1_  (.A(\v0/z1/z2/z2/temp [3]),
    .B(\v0/z1/z2/z2/temp [2]),
    .X(\v0/z1/z2/q1 [2]));
 sky130_fd_sc_hd__and2_0 \v0/z1/z2/z3/_0_  (.A(abs_b[2]),
    .B(abs_a[4]),
    .X(\v0/z1/z2/q2 [0]));
 sky130_fd_sc_hd__and2_0 \v0/z1/z2/z3/_1_  (.A(abs_b[2]),
    .B(abs_a[5]),
    .X(\v0/z1/z2/z3/temp [0]));
 sky130_fd_sc_hd__and2_0 \v0/z1/z2/z3/_2_  (.A(abs_a[4]),
    .B(abs_b[3]),
    .X(\v0/z1/z2/z3/temp [1]));
 sky130_fd_sc_hd__and2_0 \v0/z1/z2/z3/_3_  (.A(abs_a[5]),
    .B(abs_b[3]),
    .X(\v0/z1/z2/z3/temp [2]));
 sky130_fd_sc_hd__and2_0 \v0/z1/z2/z3/z1/_0_  (.A(\v0/z1/z2/z3/temp [1]),
    .B(\v0/z1/z2/z3/temp [0]),
    .X(\v0/z1/z2/z3/temp [3]));
 sky130_fd_sc_hd__xor2_1 \v0/z1/z2/z3/z1/_1_  (.A(\v0/z1/z2/z3/temp [1]),
    .B(\v0/z1/z2/z3/temp [0]),
    .X(\v0/z1/z2/q2 [1]));
 sky130_fd_sc_hd__and2_0 \v0/z1/z2/z3/z2/_0_  (.A(\v0/z1/z2/z3/temp [3]),
    .B(\v0/z1/z2/z3/temp [2]),
    .X(\v0/z1/z2/q2 [3]));
 sky130_fd_sc_hd__xor2_1 \v0/z1/z2/z3/z2/_1_  (.A(\v0/z1/z2/z3/temp [3]),
    .B(\v0/z1/z2/z3/temp [2]),
    .X(\v0/z1/z2/q2 [2]));
 sky130_fd_sc_hd__and2_0 \v0/z1/z2/z4/_0_  (.A(abs_b[2]),
    .B(abs_a[6]),
    .X(\v0/z1/z2/q3 [0]));
 sky130_fd_sc_hd__and2_0 \v0/z1/z2/z4/_1_  (.A(abs_b[2]),
    .B(abs_a[7]),
    .X(\v0/z1/z2/z4/temp [0]));
 sky130_fd_sc_hd__and2_0 \v0/z1/z2/z4/_2_  (.A(abs_a[6]),
    .B(abs_b[3]),
    .X(\v0/z1/z2/z4/temp [1]));
 sky130_fd_sc_hd__and2_0 \v0/z1/z2/z4/_3_  (.A(abs_a[7]),
    .B(abs_b[3]),
    .X(\v0/z1/z2/z4/temp [2]));
 sky130_fd_sc_hd__and2_0 \v0/z1/z2/z4/z1/_0_  (.A(\v0/z1/z2/z4/temp [1]),
    .B(\v0/z1/z2/z4/temp [0]),
    .X(\v0/z1/z2/z4/temp [3]));
 sky130_fd_sc_hd__xor2_1 \v0/z1/z2/z4/z1/_1_  (.A(\v0/z1/z2/z4/temp [1]),
    .B(\v0/z1/z2/z4/temp [0]),
    .X(\v0/z1/z2/q3 [1]));
 sky130_fd_sc_hd__and2_0 \v0/z1/z2/z4/z2/_0_  (.A(\v0/z1/z2/z4/temp [3]),
    .B(\v0/z1/z2/z4/temp [2]),
    .X(\v0/z1/z2/q3 [3]));
 sky130_fd_sc_hd__xor2_1 \v0/z1/z2/z4/z2/_1_  (.A(\v0/z1/z2/z4/temp [3]),
    .B(\v0/z1/z2/z4/temp [2]),
    .X(\v0/z1/z2/q3 [2]));
 sky130_fd_sc_hd__xnor2_1 \v0/z1/z2/z5/_07_  (.A(\v0/z1/z2/q0 [2]),
    .B(\v0/z1/z2/q1 [0]),
    .Y(\v0/z1/z2/z5/_00_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z1/z2/z5/_08_  (.A(\v0/z1/z2/_02_ ),
    .B(\v0/z1/z2/z5/_00_ ),
    .Y(\v0/z1/z2/q4 [0]));
 sky130_fd_sc_hd__maj3_1 \v0/z1/z2/z5/_09_  (.A(\v0/z1/z2/q0 [2]),
    .B(\v0/z1/z2/q1 [0]),
    .C(\v0/z1/z2/_02_ ),
    .X(\v0/z1/z2/z5/_01_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z1/z2/z5/_10_  (.A(\v0/z1/z2/q0 [3]),
    .B(\v0/z1/z2/q1 [1]),
    .Y(\v0/z1/z2/z5/_02_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z1/z2/z5/_11_  (.A(\v0/z1/z2/z5/_01_ ),
    .B(\v0/z1/z2/z5/_02_ ),
    .Y(\v0/z1/z2/q4 [1]));
 sky130_fd_sc_hd__maj3_1 \v0/z1/z2/z5/_12_  (.A(\v0/z1/z2/q0 [3]),
    .B(\v0/z1/z2/q1 [1]),
    .C(\v0/z1/z2/z5/_01_ ),
    .X(\v0/z1/z2/z5/_03_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z1/z2/z5/_13_  (.A(\v0/z1/z2/_00_ ),
    .B(\v0/z1/z2/q1 [2]),
    .Y(\v0/z1/z2/z5/_04_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z1/z2/z5/_14_  (.A(\v0/z1/z2/z5/_03_ ),
    .B(\v0/z1/z2/z5/_04_ ),
    .Y(\v0/z1/z2/q4 [2]));
 sky130_fd_sc_hd__maj3_1 \v0/z1/z2/z5/_15_  (.A(\v0/z1/z2/_00_ ),
    .B(\v0/z1/z2/q1 [2]),
    .C(\v0/z1/z2/z5/_03_ ),
    .X(\v0/z1/z2/z5/_05_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z1/z2/z5/_16_  (.A(\v0/z1/z2/_01_ ),
    .B(\v0/z1/z2/q1 [3]),
    .Y(\v0/z1/z2/z5/_06_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z1/z2/z5/_17_  (.A(\v0/z1/z2/z5/_05_ ),
    .B(\v0/z1/z2/z5/_06_ ),
    .Y(\v0/z1/z2/q4 [3]));
 sky130_fd_sc_hd__maj3_1 \v0/z1/z2/z5/_18_  (.A(\v0/z1/z2/_01_ ),
    .B(\v0/z1/z2/q1 [3]),
    .C(\v0/z1/z2/z5/_05_ ),
    .X(\v0/z1/z2/z5/Cout ));
 sky130_fd_sc_hd__xnor2_1 \v0/z1/z2/z6/_19_  (.A(\v0/z1/z2/_05_ ),
    .B(\v0/z1/z2/q2 [0]),
    .Y(\v0/z1/z2/z6/_00_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z1/z2/z6/_20_  (.A(\v0/z1/z2/_07_ ),
    .B(\v0/z1/z2/z6/_00_ ),
    .Y(\v0/z1/z2/q5 [0]));
 sky130_fd_sc_hd__maj3_1 \v0/z1/z2/z6/_21_  (.A(\v0/z1/z2/_05_ ),
    .B(\v0/z1/z2/q2 [0]),
    .C(\v0/z1/z2/_07_ ),
    .X(\v0/z1/z2/z6/_01_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z1/z2/z6/_22_  (.A(\v0/z1/z2/_06_ ),
    .B(\v0/z1/z2/q2 [1]),
    .Y(\v0/z1/z2/z6/_02_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z1/z2/z6/_23_  (.A(\v0/z1/z2/z6/_01_ ),
    .B(\v0/z1/z2/z6/_02_ ),
    .Y(\v0/z1/z2/q5 [1]));
 sky130_fd_sc_hd__maj3_1 \v0/z1/z2/z6/_24_  (.A(\v0/z1/z2/_06_ ),
    .B(\v0/z1/z2/q2 [1]),
    .C(\v0/z1/z2/z6/_01_ ),
    .X(\v0/z1/z2/z6/_03_ ));
 sky130_fd_sc_hd__lpflow_inputiso1p_1 \v0/z1/z2/z6/_25_  (.A(\v0/z1/z2/q3 [0]),
    .SLEEP(\v0/z1/z2/q2 [2]),
    .X(\v0/z1/z2/z6/_04_ ));
 sky130_fd_sc_hd__and2_0 \v0/z1/z2/z6/_26_  (.A(\v0/z1/z2/q3 [0]),
    .B(\v0/z1/z2/q2 [2]),
    .X(\v0/z1/z2/z6/_05_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z1/z2/z6/_27_  (.A(\v0/z1/z2/q3 [0]),
    .B(\v0/z1/z2/q2 [2]),
    .Y(\v0/z1/z2/z6/_06_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z1/z2/z6/_28_  (.A(\v0/z1/z2/z6/_04_ ),
    .B(\v0/z1/z2/z6/_06_ ),
    .Y(\v0/z1/z2/z6/_07_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z1/z2/z6/_29_  (.A(\v0/z1/z2/z6/_03_ ),
    .B(\v0/z1/z2/z6/_07_ ),
    .Y(\v0/z1/z2/q5 [2]));
 sky130_fd_sc_hd__nand2_1 \v0/z1/z2/z6/_30_  (.A(\v0/z1/z2/q3 [1]),
    .B(\v0/z1/z2/q2 [3]),
    .Y(\v0/z1/z2/z6/_08_ ));
 sky130_fd_sc_hd__xor2_1 \v0/z1/z2/z6/_31_  (.A(\v0/z1/z2/q3 [1]),
    .B(\v0/z1/z2/q2 [3]),
    .X(\v0/z1/z2/z6/_09_ ));
 sky130_fd_sc_hd__o21ai_0 \v0/z1/z2/z6/_32_  (.A1(\v0/z1/z2/z6/_03_ ),
    .A2(\v0/z1/z2/z6/_05_ ),
    .B1(\v0/z1/z2/z6/_04_ ),
    .Y(\v0/z1/z2/z6/_10_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z1/z2/z6/_33_  (.A(\v0/z1/z2/z6/_09_ ),
    .B(\v0/z1/z2/z6/_10_ ),
    .Y(\v0/z1/z2/q5 [3]));
 sky130_fd_sc_hd__nor2_1 \v0/z1/z2/z6/_34_  (.A(\v0/z1/z2/q3 [2]),
    .B(\v0/z1/z2/_03_ ),
    .Y(\v0/z1/z2/z6/_11_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z1/z2/z6/_35_  (.A(\v0/z1/z2/q3 [2]),
    .B(\v0/z1/z2/_03_ ),
    .Y(\v0/z1/z2/z6/_12_ ));
 sky130_fd_sc_hd__nand2b_1 \v0/z1/z2/z6/_36_  (.A_N(\v0/z1/z2/z6/_11_ ),
    .B(\v0/z1/z2/z6/_12_ ),
    .Y(\v0/z1/z2/z6/_13_ ));
 sky130_fd_sc_hd__o221ai_1 \v0/z1/z2/z6/_37_  (.A1(\v0/z1/z2/q3 [1]),
    .A2(\v0/z1/z2/q2 [3]),
    .B1(\v0/z1/z2/z6/_03_ ),
    .B2(\v0/z1/z2/z6/_05_ ),
    .C1(\v0/z1/z2/z6/_04_ ),
    .Y(\v0/z1/z2/z6/_14_ ));
 sky130_fd_sc_hd__a21oi_1 \v0/z1/z2/z6/_38_  (.A1(\v0/z1/z2/z6/_08_ ),
    .A2(\v0/z1/z2/z6/_14_ ),
    .B1(\v0/z1/z2/z6/_13_ ),
    .Y(\v0/z1/z2/z6/_15_ ));
 sky130_fd_sc_hd__and3_1 \v0/z1/z2/z6/_39_  (.A(\v0/z1/z2/z6/_08_ ),
    .B(\v0/z1/z2/z6/_13_ ),
    .C(\v0/z1/z2/z6/_14_ ),
    .X(\v0/z1/z2/z6/_16_ ));
 sky130_fd_sc_hd__nor2_1 \v0/z1/z2/z6/_40_  (.A(\v0/z1/z2/z6/_15_ ),
    .B(\v0/z1/z2/z6/_16_ ),
    .Y(\v0/z1/z2/q5 [4]));
 sky130_fd_sc_hd__xnor2_1 \v0/z1/z2/z6/_41_  (.A(\v0/z1/z2/q3 [3]),
    .B(\v0/z1/z2/_04_ ),
    .Y(\v0/z1/z2/z6/_17_ ));
 sky130_fd_sc_hd__a31oi_1 \v0/z1/z2/z6/_42_  (.A1(\v0/z1/z2/z6/_08_ ),
    .A2(\v0/z1/z2/z6/_12_ ),
    .A3(\v0/z1/z2/z6/_14_ ),
    .B1(\v0/z1/z2/z6/_11_ ),
    .Y(\v0/z1/z2/z6/_18_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z1/z2/z6/_43_  (.A(\v0/z1/z2/z6/_17_ ),
    .B(\v0/z1/z2/z6/_18_ ),
    .Y(\v0/z1/z2/q5 [5]));
 sky130_fd_sc_hd__maj3_1 \v0/z1/z2/z6/_44_  (.A(\v0/z1/z2/q3 [3]),
    .B(\v0/z1/z2/_04_ ),
    .C(\v0/z1/z2/z6/_18_ ),
    .X(\v0/z1/z2/z6/Cout ));
 sky130_fd_sc_hd__xnor2_1 \v0/z1/z2/z7/_19_  (.A(\v0/z1/z2/q5 [0]),
    .B(\v0/z1/z2/q4 [0]),
    .Y(\v0/z1/z2/z7/_00_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z1/z2/z7/_20_  (.A(\v0/z1/z2/_10_ ),
    .B(\v0/z1/z2/z7/_00_ ),
    .Y(\v0/z1/q1 [2]));
 sky130_fd_sc_hd__maj3_1 \v0/z1/z2/z7/_21_  (.A(\v0/z1/z2/q5 [0]),
    .B(\v0/z1/z2/q4 [0]),
    .C(\v0/z1/z2/_10_ ),
    .X(\v0/z1/z2/z7/_01_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z1/z2/z7/_22_  (.A(\v0/z1/z2/q5 [1]),
    .B(\v0/z1/z2/q4 [1]),
    .Y(\v0/z1/z2/z7/_02_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z1/z2/z7/_23_  (.A(\v0/z1/z2/z7/_01_ ),
    .B(\v0/z1/z2/z7/_02_ ),
    .Y(\v0/z1/q1 [3]));
 sky130_fd_sc_hd__maj3_1 \v0/z1/z2/z7/_24_  (.A(\v0/z1/z2/q5 [1]),
    .B(\v0/z1/z2/q4 [1]),
    .C(\v0/z1/z2/z7/_01_ ),
    .X(\v0/z1/z2/z7/_03_ ));
 sky130_fd_sc_hd__lpflow_inputiso1p_1 \v0/z1/z2/z7/_25_  (.A(\v0/z1/z2/q5 [2]),
    .SLEEP(\v0/z1/z2/q4 [2]),
    .X(\v0/z1/z2/z7/_04_ ));
 sky130_fd_sc_hd__and2_0 \v0/z1/z2/z7/_26_  (.A(\v0/z1/z2/q5 [2]),
    .B(\v0/z1/z2/q4 [2]),
    .X(\v0/z1/z2/z7/_05_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z1/z2/z7/_27_  (.A(\v0/z1/z2/q5 [2]),
    .B(\v0/z1/z2/q4 [2]),
    .Y(\v0/z1/z2/z7/_06_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z1/z2/z7/_28_  (.A(\v0/z1/z2/z7/_04_ ),
    .B(\v0/z1/z2/z7/_06_ ),
    .Y(\v0/z1/z2/z7/_07_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z1/z2/z7/_29_  (.A(\v0/z1/z2/z7/_03_ ),
    .B(\v0/z1/z2/z7/_07_ ),
    .Y(\v0/z1/q1 [4]));
 sky130_fd_sc_hd__nand2_1 \v0/z1/z2/z7/_30_  (.A(\v0/z1/z2/q5 [3]),
    .B(\v0/z1/z2/q4 [3]),
    .Y(\v0/z1/z2/z7/_08_ ));
 sky130_fd_sc_hd__xor2_1 \v0/z1/z2/z7/_31_  (.A(\v0/z1/z2/q5 [3]),
    .B(\v0/z1/z2/q4 [3]),
    .X(\v0/z1/z2/z7/_09_ ));
 sky130_fd_sc_hd__o21ai_0 \v0/z1/z2/z7/_32_  (.A1(\v0/z1/z2/z7/_03_ ),
    .A2(\v0/z1/z2/z7/_05_ ),
    .B1(\v0/z1/z2/z7/_04_ ),
    .Y(\v0/z1/z2/z7/_10_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z1/z2/z7/_33_  (.A(\v0/z1/z2/z7/_09_ ),
    .B(\v0/z1/z2/z7/_10_ ),
    .Y(\v0/z1/q1 [5]));
 sky130_fd_sc_hd__nor2_1 \v0/z1/z2/z7/_34_  (.A(\v0/z1/z2/q5 [4]),
    .B(\v0/z1/z2/_08_ ),
    .Y(\v0/z1/z2/z7/_11_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z1/z2/z7/_35_  (.A(\v0/z1/z2/q5 [4]),
    .B(\v0/z1/z2/_08_ ),
    .Y(\v0/z1/z2/z7/_12_ ));
 sky130_fd_sc_hd__nand2b_1 \v0/z1/z2/z7/_36_  (.A_N(\v0/z1/z2/z7/_11_ ),
    .B(\v0/z1/z2/z7/_12_ ),
    .Y(\v0/z1/z2/z7/_13_ ));
 sky130_fd_sc_hd__o221ai_1 \v0/z1/z2/z7/_37_  (.A1(\v0/z1/z2/q5 [3]),
    .A2(\v0/z1/z2/q4 [3]),
    .B1(\v0/z1/z2/z7/_03_ ),
    .B2(\v0/z1/z2/z7/_05_ ),
    .C1(\v0/z1/z2/z7/_04_ ),
    .Y(\v0/z1/z2/z7/_14_ ));
 sky130_fd_sc_hd__a21oi_1 \v0/z1/z2/z7/_38_  (.A1(\v0/z1/z2/z7/_08_ ),
    .A2(\v0/z1/z2/z7/_14_ ),
    .B1(\v0/z1/z2/z7/_13_ ),
    .Y(\v0/z1/z2/z7/_15_ ));
 sky130_fd_sc_hd__and3_1 \v0/z1/z2/z7/_39_  (.A(\v0/z1/z2/z7/_08_ ),
    .B(\v0/z1/z2/z7/_13_ ),
    .C(\v0/z1/z2/z7/_14_ ),
    .X(\v0/z1/z2/z7/_16_ ));
 sky130_fd_sc_hd__nor2_1 \v0/z1/z2/z7/_40_  (.A(\v0/z1/z2/z7/_15_ ),
    .B(\v0/z1/z2/z7/_16_ ),
    .Y(\v0/z1/q1 [6]));
 sky130_fd_sc_hd__xnor2_1 \v0/z1/z2/z7/_41_  (.A(\v0/z1/z2/q5 [5]),
    .B(\v0/z1/z2/_09_ ),
    .Y(\v0/z1/z2/z7/_17_ ));
 sky130_fd_sc_hd__a31oi_1 \v0/z1/z2/z7/_42_  (.A1(\v0/z1/z2/z7/_08_ ),
    .A2(\v0/z1/z2/z7/_12_ ),
    .A3(\v0/z1/z2/z7/_14_ ),
    .B1(\v0/z1/z2/z7/_11_ ),
    .Y(\v0/z1/z2/z7/_18_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z1/z2/z7/_43_  (.A(\v0/z1/z2/z7/_17_ ),
    .B(\v0/z1/z2/z7/_18_ ),
    .Y(\v0/z1/q1 [7]));
 sky130_fd_sc_hd__maj3_1 \v0/z1/z2/z7/_44_  (.A(\v0/z1/z2/q5 [5]),
    .B(\v0/z1/z2/_09_ ),
    .C(\v0/z1/z2/z7/_18_ ),
    .X(\v0/z1/z2/z7/Cout ));
 sky130_fd_sc_hd__conb_1 \v0/z1/z3/_11_  (.LO(\v0/z1/z3/_00_ ));
 sky130_fd_sc_hd__conb_1 \v0/z1/z3/_12_  (.LO(\v0/z1/z3/_01_ ));
 sky130_fd_sc_hd__conb_1 \v0/z1/z3/_13_  (.LO(\v0/z1/z3/_02_ ));
 sky130_fd_sc_hd__conb_1 \v0/z1/z3/_14_  (.LO(\v0/z1/z3/_03_ ));
 sky130_fd_sc_hd__conb_1 \v0/z1/z3/_15_  (.LO(\v0/z1/z3/_04_ ));
 sky130_fd_sc_hd__conb_1 \v0/z1/z3/_16_  (.LO(\v0/z1/z3/_05_ ));
 sky130_fd_sc_hd__conb_1 \v0/z1/z3/_17_  (.LO(\v0/z1/z3/_06_ ));
 sky130_fd_sc_hd__conb_1 \v0/z1/z3/_18_  (.LO(\v0/z1/z3/_07_ ));
 sky130_fd_sc_hd__conb_1 \v0/z1/z3/_19_  (.LO(\v0/z1/z3/_08_ ));
 sky130_fd_sc_hd__conb_1 \v0/z1/z3/_20_  (.LO(\v0/z1/z3/_09_ ));
 sky130_fd_sc_hd__conb_1 \v0/z1/z3/_21_  (.LO(\v0/z1/z3/_10_ ));
 sky130_fd_sc_hd__and2_0 \v0/z1/z3/z1/_0_  (.A(abs_b[4]),
    .B(a[0]),
    .X(\v0/z1/q2 [0]));
 sky130_fd_sc_hd__and2_0 \v0/z1/z3/z1/_1_  (.A(abs_b[4]),
    .B(abs_a[1]),
    .X(\v0/z1/z3/z1/temp [0]));
 sky130_fd_sc_hd__and2_0 \v0/z1/z3/z1/_2_  (.A(a[0]),
    .B(abs_b[5]),
    .X(\v0/z1/z3/z1/temp [1]));
 sky130_fd_sc_hd__and2_0 \v0/z1/z3/z1/_3_  (.A(abs_a[1]),
    .B(abs_b[5]),
    .X(\v0/z1/z3/z1/temp [2]));
 sky130_fd_sc_hd__and2_0 \v0/z1/z3/z1/z1/_0_  (.A(\v0/z1/z3/z1/temp [1]),
    .B(\v0/z1/z3/z1/temp [0]),
    .X(\v0/z1/z3/z1/temp [3]));
 sky130_fd_sc_hd__xor2_1 \v0/z1/z3/z1/z1/_1_  (.A(\v0/z1/z3/z1/temp [1]),
    .B(\v0/z1/z3/z1/temp [0]),
    .X(\v0/z1/q2 [1]));
 sky130_fd_sc_hd__and2_0 \v0/z1/z3/z1/z2/_0_  (.A(\v0/z1/z3/z1/temp [3]),
    .B(\v0/z1/z3/z1/temp [2]),
    .X(\v0/z1/z3/q0 [3]));
 sky130_fd_sc_hd__xor2_1 \v0/z1/z3/z1/z2/_1_  (.A(\v0/z1/z3/z1/temp [3]),
    .B(\v0/z1/z3/z1/temp [2]),
    .X(\v0/z1/z3/q0 [2]));
 sky130_fd_sc_hd__and2_0 \v0/z1/z3/z2/_0_  (.A(abs_b[4]),
    .B(abs_a[2]),
    .X(\v0/z1/z3/q1 [0]));
 sky130_fd_sc_hd__and2_0 \v0/z1/z3/z2/_1_  (.A(abs_b[4]),
    .B(abs_a[3]),
    .X(\v0/z1/z3/z2/temp [0]));
 sky130_fd_sc_hd__and2_0 \v0/z1/z3/z2/_2_  (.A(abs_a[2]),
    .B(abs_b[5]),
    .X(\v0/z1/z3/z2/temp [1]));
 sky130_fd_sc_hd__and2_0 \v0/z1/z3/z2/_3_  (.A(abs_a[3]),
    .B(abs_b[5]),
    .X(\v0/z1/z3/z2/temp [2]));
 sky130_fd_sc_hd__and2_0 \v0/z1/z3/z2/z1/_0_  (.A(\v0/z1/z3/z2/temp [1]),
    .B(\v0/z1/z3/z2/temp [0]),
    .X(\v0/z1/z3/z2/temp [3]));
 sky130_fd_sc_hd__xor2_1 \v0/z1/z3/z2/z1/_1_  (.A(\v0/z1/z3/z2/temp [1]),
    .B(\v0/z1/z3/z2/temp [0]),
    .X(\v0/z1/z3/q1 [1]));
 sky130_fd_sc_hd__and2_0 \v0/z1/z3/z2/z2/_0_  (.A(\v0/z1/z3/z2/temp [3]),
    .B(\v0/z1/z3/z2/temp [2]),
    .X(\v0/z1/z3/q1 [3]));
 sky130_fd_sc_hd__xor2_1 \v0/z1/z3/z2/z2/_1_  (.A(\v0/z1/z3/z2/temp [3]),
    .B(\v0/z1/z3/z2/temp [2]),
    .X(\v0/z1/z3/q1 [2]));
 sky130_fd_sc_hd__and2_0 \v0/z1/z3/z3/_0_  (.A(abs_b[6]),
    .B(a[0]),
    .X(\v0/z1/z3/q2 [0]));
 sky130_fd_sc_hd__and2_0 \v0/z1/z3/z3/_1_  (.A(abs_b[6]),
    .B(abs_a[1]),
    .X(\v0/z1/z3/z3/temp [0]));
 sky130_fd_sc_hd__and2_0 \v0/z1/z3/z3/_2_  (.A(a[0]),
    .B(abs_b[7]),
    .X(\v0/z1/z3/z3/temp [1]));
 sky130_fd_sc_hd__and2_0 \v0/z1/z3/z3/_3_  (.A(abs_a[1]),
    .B(abs_b[7]),
    .X(\v0/z1/z3/z3/temp [2]));
 sky130_fd_sc_hd__and2_0 \v0/z1/z3/z3/z1/_0_  (.A(\v0/z1/z3/z3/temp [1]),
    .B(\v0/z1/z3/z3/temp [0]),
    .X(\v0/z1/z3/z3/temp [3]));
 sky130_fd_sc_hd__xor2_1 \v0/z1/z3/z3/z1/_1_  (.A(\v0/z1/z3/z3/temp [1]),
    .B(\v0/z1/z3/z3/temp [0]),
    .X(\v0/z1/z3/q2 [1]));
 sky130_fd_sc_hd__and2_0 \v0/z1/z3/z3/z2/_0_  (.A(\v0/z1/z3/z3/temp [3]),
    .B(\v0/z1/z3/z3/temp [2]),
    .X(\v0/z1/z3/q2 [3]));
 sky130_fd_sc_hd__xor2_1 \v0/z1/z3/z3/z2/_1_  (.A(\v0/z1/z3/z3/temp [3]),
    .B(\v0/z1/z3/z3/temp [2]),
    .X(\v0/z1/z3/q2 [2]));
 sky130_fd_sc_hd__and2_0 \v0/z1/z3/z4/_0_  (.A(abs_b[6]),
    .B(abs_a[2]),
    .X(\v0/z1/z3/q3 [0]));
 sky130_fd_sc_hd__and2_0 \v0/z1/z3/z4/_1_  (.A(abs_b[6]),
    .B(abs_a[3]),
    .X(\v0/z1/z3/z4/temp [0]));
 sky130_fd_sc_hd__and2_0 \v0/z1/z3/z4/_2_  (.A(abs_a[2]),
    .B(abs_b[7]),
    .X(\v0/z1/z3/z4/temp [1]));
 sky130_fd_sc_hd__and2_0 \v0/z1/z3/z4/_3_  (.A(abs_a[3]),
    .B(abs_b[7]),
    .X(\v0/z1/z3/z4/temp [2]));
 sky130_fd_sc_hd__and2_0 \v0/z1/z3/z4/z1/_0_  (.A(\v0/z1/z3/z4/temp [1]),
    .B(\v0/z1/z3/z4/temp [0]),
    .X(\v0/z1/z3/z4/temp [3]));
 sky130_fd_sc_hd__xor2_1 \v0/z1/z3/z4/z1/_1_  (.A(\v0/z1/z3/z4/temp [1]),
    .B(\v0/z1/z3/z4/temp [0]),
    .X(\v0/z1/z3/q3 [1]));
 sky130_fd_sc_hd__and2_0 \v0/z1/z3/z4/z2/_0_  (.A(\v0/z1/z3/z4/temp [3]),
    .B(\v0/z1/z3/z4/temp [2]),
    .X(\v0/z1/z3/q3 [3]));
 sky130_fd_sc_hd__xor2_1 \v0/z1/z3/z4/z2/_1_  (.A(\v0/z1/z3/z4/temp [3]),
    .B(\v0/z1/z3/z4/temp [2]),
    .X(\v0/z1/z3/q3 [2]));
 sky130_fd_sc_hd__xnor2_1 \v0/z1/z3/z5/_07_  (.A(\v0/z1/z3/q0 [2]),
    .B(\v0/z1/z3/q1 [0]),
    .Y(\v0/z1/z3/z5/_00_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z1/z3/z5/_08_  (.A(\v0/z1/z3/_02_ ),
    .B(\v0/z1/z3/z5/_00_ ),
    .Y(\v0/z1/z3/q4 [0]));
 sky130_fd_sc_hd__maj3_1 \v0/z1/z3/z5/_09_  (.A(\v0/z1/z3/q0 [2]),
    .B(\v0/z1/z3/q1 [0]),
    .C(\v0/z1/z3/_02_ ),
    .X(\v0/z1/z3/z5/_01_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z1/z3/z5/_10_  (.A(\v0/z1/z3/q0 [3]),
    .B(\v0/z1/z3/q1 [1]),
    .Y(\v0/z1/z3/z5/_02_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z1/z3/z5/_11_  (.A(\v0/z1/z3/z5/_01_ ),
    .B(\v0/z1/z3/z5/_02_ ),
    .Y(\v0/z1/z3/q4 [1]));
 sky130_fd_sc_hd__maj3_1 \v0/z1/z3/z5/_12_  (.A(\v0/z1/z3/q0 [3]),
    .B(\v0/z1/z3/q1 [1]),
    .C(\v0/z1/z3/z5/_01_ ),
    .X(\v0/z1/z3/z5/_03_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z1/z3/z5/_13_  (.A(\v0/z1/z3/_00_ ),
    .B(\v0/z1/z3/q1 [2]),
    .Y(\v0/z1/z3/z5/_04_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z1/z3/z5/_14_  (.A(\v0/z1/z3/z5/_03_ ),
    .B(\v0/z1/z3/z5/_04_ ),
    .Y(\v0/z1/z3/q4 [2]));
 sky130_fd_sc_hd__maj3_1 \v0/z1/z3/z5/_15_  (.A(\v0/z1/z3/_00_ ),
    .B(\v0/z1/z3/q1 [2]),
    .C(\v0/z1/z3/z5/_03_ ),
    .X(\v0/z1/z3/z5/_05_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z1/z3/z5/_16_  (.A(\v0/z1/z3/_01_ ),
    .B(\v0/z1/z3/q1 [3]),
    .Y(\v0/z1/z3/z5/_06_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z1/z3/z5/_17_  (.A(\v0/z1/z3/z5/_05_ ),
    .B(\v0/z1/z3/z5/_06_ ),
    .Y(\v0/z1/z3/q4 [3]));
 sky130_fd_sc_hd__maj3_1 \v0/z1/z3/z5/_18_  (.A(\v0/z1/z3/_01_ ),
    .B(\v0/z1/z3/q1 [3]),
    .C(\v0/z1/z3/z5/_05_ ),
    .X(\v0/z1/z3/z5/Cout ));
 sky130_fd_sc_hd__xnor2_1 \v0/z1/z3/z6/_19_  (.A(\v0/z1/z3/_05_ ),
    .B(\v0/z1/z3/q2 [0]),
    .Y(\v0/z1/z3/z6/_00_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z1/z3/z6/_20_  (.A(\v0/z1/z3/_07_ ),
    .B(\v0/z1/z3/z6/_00_ ),
    .Y(\v0/z1/z3/q5 [0]));
 sky130_fd_sc_hd__maj3_1 \v0/z1/z3/z6/_21_  (.A(\v0/z1/z3/_05_ ),
    .B(\v0/z1/z3/q2 [0]),
    .C(\v0/z1/z3/_07_ ),
    .X(\v0/z1/z3/z6/_01_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z1/z3/z6/_22_  (.A(\v0/z1/z3/_06_ ),
    .B(\v0/z1/z3/q2 [1]),
    .Y(\v0/z1/z3/z6/_02_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z1/z3/z6/_23_  (.A(\v0/z1/z3/z6/_01_ ),
    .B(\v0/z1/z3/z6/_02_ ),
    .Y(\v0/z1/z3/q5 [1]));
 sky130_fd_sc_hd__maj3_1 \v0/z1/z3/z6/_24_  (.A(\v0/z1/z3/_06_ ),
    .B(\v0/z1/z3/q2 [1]),
    .C(\v0/z1/z3/z6/_01_ ),
    .X(\v0/z1/z3/z6/_03_ ));
 sky130_fd_sc_hd__lpflow_inputiso1p_1 \v0/z1/z3/z6/_25_  (.A(\v0/z1/z3/q3 [0]),
    .SLEEP(\v0/z1/z3/q2 [2]),
    .X(\v0/z1/z3/z6/_04_ ));
 sky130_fd_sc_hd__and2_0 \v0/z1/z3/z6/_26_  (.A(\v0/z1/z3/q3 [0]),
    .B(\v0/z1/z3/q2 [2]),
    .X(\v0/z1/z3/z6/_05_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z1/z3/z6/_27_  (.A(\v0/z1/z3/q3 [0]),
    .B(\v0/z1/z3/q2 [2]),
    .Y(\v0/z1/z3/z6/_06_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z1/z3/z6/_28_  (.A(\v0/z1/z3/z6/_04_ ),
    .B(\v0/z1/z3/z6/_06_ ),
    .Y(\v0/z1/z3/z6/_07_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z1/z3/z6/_29_  (.A(\v0/z1/z3/z6/_03_ ),
    .B(\v0/z1/z3/z6/_07_ ),
    .Y(\v0/z1/z3/q5 [2]));
 sky130_fd_sc_hd__nand2_1 \v0/z1/z3/z6/_30_  (.A(\v0/z1/z3/q3 [1]),
    .B(\v0/z1/z3/q2 [3]),
    .Y(\v0/z1/z3/z6/_08_ ));
 sky130_fd_sc_hd__xor2_1 \v0/z1/z3/z6/_31_  (.A(\v0/z1/z3/q3 [1]),
    .B(\v0/z1/z3/q2 [3]),
    .X(\v0/z1/z3/z6/_09_ ));
 sky130_fd_sc_hd__o21ai_0 \v0/z1/z3/z6/_32_  (.A1(\v0/z1/z3/z6/_03_ ),
    .A2(\v0/z1/z3/z6/_05_ ),
    .B1(\v0/z1/z3/z6/_04_ ),
    .Y(\v0/z1/z3/z6/_10_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z1/z3/z6/_33_  (.A(\v0/z1/z3/z6/_09_ ),
    .B(\v0/z1/z3/z6/_10_ ),
    .Y(\v0/z1/z3/q5 [3]));
 sky130_fd_sc_hd__nor2_1 \v0/z1/z3/z6/_34_  (.A(\v0/z1/z3/q3 [2]),
    .B(\v0/z1/z3/_03_ ),
    .Y(\v0/z1/z3/z6/_11_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z1/z3/z6/_35_  (.A(\v0/z1/z3/q3 [2]),
    .B(\v0/z1/z3/_03_ ),
    .Y(\v0/z1/z3/z6/_12_ ));
 sky130_fd_sc_hd__nand2b_1 \v0/z1/z3/z6/_36_  (.A_N(\v0/z1/z3/z6/_11_ ),
    .B(\v0/z1/z3/z6/_12_ ),
    .Y(\v0/z1/z3/z6/_13_ ));
 sky130_fd_sc_hd__o221ai_1 \v0/z1/z3/z6/_37_  (.A1(\v0/z1/z3/q3 [1]),
    .A2(\v0/z1/z3/q2 [3]),
    .B1(\v0/z1/z3/z6/_03_ ),
    .B2(\v0/z1/z3/z6/_05_ ),
    .C1(\v0/z1/z3/z6/_04_ ),
    .Y(\v0/z1/z3/z6/_14_ ));
 sky130_fd_sc_hd__a21oi_1 \v0/z1/z3/z6/_38_  (.A1(\v0/z1/z3/z6/_08_ ),
    .A2(\v0/z1/z3/z6/_14_ ),
    .B1(\v0/z1/z3/z6/_13_ ),
    .Y(\v0/z1/z3/z6/_15_ ));
 sky130_fd_sc_hd__and3_1 \v0/z1/z3/z6/_39_  (.A(\v0/z1/z3/z6/_08_ ),
    .B(\v0/z1/z3/z6/_13_ ),
    .C(\v0/z1/z3/z6/_14_ ),
    .X(\v0/z1/z3/z6/_16_ ));
 sky130_fd_sc_hd__nor2_1 \v0/z1/z3/z6/_40_  (.A(\v0/z1/z3/z6/_15_ ),
    .B(\v0/z1/z3/z6/_16_ ),
    .Y(\v0/z1/z3/q5 [4]));
 sky130_fd_sc_hd__xnor2_1 \v0/z1/z3/z6/_41_  (.A(\v0/z1/z3/q3 [3]),
    .B(\v0/z1/z3/_04_ ),
    .Y(\v0/z1/z3/z6/_17_ ));
 sky130_fd_sc_hd__a31oi_1 \v0/z1/z3/z6/_42_  (.A1(\v0/z1/z3/z6/_08_ ),
    .A2(\v0/z1/z3/z6/_12_ ),
    .A3(\v0/z1/z3/z6/_14_ ),
    .B1(\v0/z1/z3/z6/_11_ ),
    .Y(\v0/z1/z3/z6/_18_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z1/z3/z6/_43_  (.A(\v0/z1/z3/z6/_17_ ),
    .B(\v0/z1/z3/z6/_18_ ),
    .Y(\v0/z1/z3/q5 [5]));
 sky130_fd_sc_hd__maj3_1 \v0/z1/z3/z6/_44_  (.A(\v0/z1/z3/q3 [3]),
    .B(\v0/z1/z3/_04_ ),
    .C(\v0/z1/z3/z6/_18_ ),
    .X(\v0/z1/z3/z6/Cout ));
 sky130_fd_sc_hd__xnor2_1 \v0/z1/z3/z7/_19_  (.A(\v0/z1/z3/q5 [0]),
    .B(\v0/z1/z3/q4 [0]),
    .Y(\v0/z1/z3/z7/_00_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z1/z3/z7/_20_  (.A(\v0/z1/z3/_10_ ),
    .B(\v0/z1/z3/z7/_00_ ),
    .Y(\v0/z1/q2 [2]));
 sky130_fd_sc_hd__maj3_1 \v0/z1/z3/z7/_21_  (.A(\v0/z1/z3/q5 [0]),
    .B(\v0/z1/z3/q4 [0]),
    .C(\v0/z1/z3/_10_ ),
    .X(\v0/z1/z3/z7/_01_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z1/z3/z7/_22_  (.A(\v0/z1/z3/q5 [1]),
    .B(\v0/z1/z3/q4 [1]),
    .Y(\v0/z1/z3/z7/_02_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z1/z3/z7/_23_  (.A(\v0/z1/z3/z7/_01_ ),
    .B(\v0/z1/z3/z7/_02_ ),
    .Y(\v0/z1/q2 [3]));
 sky130_fd_sc_hd__maj3_1 \v0/z1/z3/z7/_24_  (.A(\v0/z1/z3/q5 [1]),
    .B(\v0/z1/z3/q4 [1]),
    .C(\v0/z1/z3/z7/_01_ ),
    .X(\v0/z1/z3/z7/_03_ ));
 sky130_fd_sc_hd__lpflow_inputiso1p_1 \v0/z1/z3/z7/_25_  (.A(\v0/z1/z3/q5 [2]),
    .SLEEP(\v0/z1/z3/q4 [2]),
    .X(\v0/z1/z3/z7/_04_ ));
 sky130_fd_sc_hd__and2_0 \v0/z1/z3/z7/_26_  (.A(\v0/z1/z3/q5 [2]),
    .B(\v0/z1/z3/q4 [2]),
    .X(\v0/z1/z3/z7/_05_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z1/z3/z7/_27_  (.A(\v0/z1/z3/q5 [2]),
    .B(\v0/z1/z3/q4 [2]),
    .Y(\v0/z1/z3/z7/_06_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z1/z3/z7/_28_  (.A(\v0/z1/z3/z7/_04_ ),
    .B(\v0/z1/z3/z7/_06_ ),
    .Y(\v0/z1/z3/z7/_07_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z1/z3/z7/_29_  (.A(\v0/z1/z3/z7/_03_ ),
    .B(\v0/z1/z3/z7/_07_ ),
    .Y(\v0/z1/q2 [4]));
 sky130_fd_sc_hd__nand2_1 \v0/z1/z3/z7/_30_  (.A(\v0/z1/z3/q5 [3]),
    .B(\v0/z1/z3/q4 [3]),
    .Y(\v0/z1/z3/z7/_08_ ));
 sky130_fd_sc_hd__xor2_1 \v0/z1/z3/z7/_31_  (.A(\v0/z1/z3/q5 [3]),
    .B(\v0/z1/z3/q4 [3]),
    .X(\v0/z1/z3/z7/_09_ ));
 sky130_fd_sc_hd__o21ai_0 \v0/z1/z3/z7/_32_  (.A1(\v0/z1/z3/z7/_03_ ),
    .A2(\v0/z1/z3/z7/_05_ ),
    .B1(\v0/z1/z3/z7/_04_ ),
    .Y(\v0/z1/z3/z7/_10_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z1/z3/z7/_33_  (.A(\v0/z1/z3/z7/_09_ ),
    .B(\v0/z1/z3/z7/_10_ ),
    .Y(\v0/z1/q2 [5]));
 sky130_fd_sc_hd__nor2_1 \v0/z1/z3/z7/_34_  (.A(\v0/z1/z3/q5 [4]),
    .B(\v0/z1/z3/_08_ ),
    .Y(\v0/z1/z3/z7/_11_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z1/z3/z7/_35_  (.A(\v0/z1/z3/q5 [4]),
    .B(\v0/z1/z3/_08_ ),
    .Y(\v0/z1/z3/z7/_12_ ));
 sky130_fd_sc_hd__nand2b_1 \v0/z1/z3/z7/_36_  (.A_N(\v0/z1/z3/z7/_11_ ),
    .B(\v0/z1/z3/z7/_12_ ),
    .Y(\v0/z1/z3/z7/_13_ ));
 sky130_fd_sc_hd__o221ai_1 \v0/z1/z3/z7/_37_  (.A1(\v0/z1/z3/q5 [3]),
    .A2(\v0/z1/z3/q4 [3]),
    .B1(\v0/z1/z3/z7/_03_ ),
    .B2(\v0/z1/z3/z7/_05_ ),
    .C1(\v0/z1/z3/z7/_04_ ),
    .Y(\v0/z1/z3/z7/_14_ ));
 sky130_fd_sc_hd__a21oi_1 \v0/z1/z3/z7/_38_  (.A1(\v0/z1/z3/z7/_08_ ),
    .A2(\v0/z1/z3/z7/_14_ ),
    .B1(\v0/z1/z3/z7/_13_ ),
    .Y(\v0/z1/z3/z7/_15_ ));
 sky130_fd_sc_hd__and3_1 \v0/z1/z3/z7/_39_  (.A(\v0/z1/z3/z7/_08_ ),
    .B(\v0/z1/z3/z7/_13_ ),
    .C(\v0/z1/z3/z7/_14_ ),
    .X(\v0/z1/z3/z7/_16_ ));
 sky130_fd_sc_hd__nor2_1 \v0/z1/z3/z7/_40_  (.A(\v0/z1/z3/z7/_15_ ),
    .B(\v0/z1/z3/z7/_16_ ),
    .Y(\v0/z1/q2 [6]));
 sky130_fd_sc_hd__xnor2_1 \v0/z1/z3/z7/_41_  (.A(\v0/z1/z3/q5 [5]),
    .B(\v0/z1/z3/_09_ ),
    .Y(\v0/z1/z3/z7/_17_ ));
 sky130_fd_sc_hd__a31oi_1 \v0/z1/z3/z7/_42_  (.A1(\v0/z1/z3/z7/_08_ ),
    .A2(\v0/z1/z3/z7/_12_ ),
    .A3(\v0/z1/z3/z7/_14_ ),
    .B1(\v0/z1/z3/z7/_11_ ),
    .Y(\v0/z1/z3/z7/_18_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z1/z3/z7/_43_  (.A(\v0/z1/z3/z7/_17_ ),
    .B(\v0/z1/z3/z7/_18_ ),
    .Y(\v0/z1/q2 [7]));
 sky130_fd_sc_hd__maj3_1 \v0/z1/z3/z7/_44_  (.A(\v0/z1/z3/q5 [5]),
    .B(\v0/z1/z3/_09_ ),
    .C(\v0/z1/z3/z7/_18_ ),
    .X(\v0/z1/z3/z7/Cout ));
 sky130_fd_sc_hd__conb_1 \v0/z1/z4/_11_  (.LO(\v0/z1/z4/_00_ ));
 sky130_fd_sc_hd__conb_1 \v0/z1/z4/_12_  (.LO(\v0/z1/z4/_01_ ));
 sky130_fd_sc_hd__conb_1 \v0/z1/z4/_13_  (.LO(\v0/z1/z4/_02_ ));
 sky130_fd_sc_hd__conb_1 \v0/z1/z4/_14_  (.LO(\v0/z1/z4/_03_ ));
 sky130_fd_sc_hd__conb_1 \v0/z1/z4/_15_  (.LO(\v0/z1/z4/_04_ ));
 sky130_fd_sc_hd__conb_1 \v0/z1/z4/_16_  (.LO(\v0/z1/z4/_05_ ));
 sky130_fd_sc_hd__conb_1 \v0/z1/z4/_17_  (.LO(\v0/z1/z4/_06_ ));
 sky130_fd_sc_hd__conb_1 \v0/z1/z4/_18_  (.LO(\v0/z1/z4/_07_ ));
 sky130_fd_sc_hd__conb_1 \v0/z1/z4/_19_  (.LO(\v0/z1/z4/_08_ ));
 sky130_fd_sc_hd__conb_1 \v0/z1/z4/_20_  (.LO(\v0/z1/z4/_09_ ));
 sky130_fd_sc_hd__conb_1 \v0/z1/z4/_21_  (.LO(\v0/z1/z4/_10_ ));
 sky130_fd_sc_hd__and2_0 \v0/z1/z4/z1/_0_  (.A(abs_b[4]),
    .B(abs_a[4]),
    .X(\v0/z1/q3 [0]));
 sky130_fd_sc_hd__and2_0 \v0/z1/z4/z1/_1_  (.A(abs_b[4]),
    .B(abs_a[5]),
    .X(\v0/z1/z4/z1/temp [0]));
 sky130_fd_sc_hd__and2_0 \v0/z1/z4/z1/_2_  (.A(abs_a[4]),
    .B(abs_b[5]),
    .X(\v0/z1/z4/z1/temp [1]));
 sky130_fd_sc_hd__and2_0 \v0/z1/z4/z1/_3_  (.A(abs_a[5]),
    .B(abs_b[5]),
    .X(\v0/z1/z4/z1/temp [2]));
 sky130_fd_sc_hd__and2_0 \v0/z1/z4/z1/z1/_0_  (.A(\v0/z1/z4/z1/temp [1]),
    .B(\v0/z1/z4/z1/temp [0]),
    .X(\v0/z1/z4/z1/temp [3]));
 sky130_fd_sc_hd__xor2_1 \v0/z1/z4/z1/z1/_1_  (.A(\v0/z1/z4/z1/temp [1]),
    .B(\v0/z1/z4/z1/temp [0]),
    .X(\v0/z1/q3 [1]));
 sky130_fd_sc_hd__and2_0 \v0/z1/z4/z1/z2/_0_  (.A(\v0/z1/z4/z1/temp [3]),
    .B(\v0/z1/z4/z1/temp [2]),
    .X(\v0/z1/z4/q0 [3]));
 sky130_fd_sc_hd__xor2_1 \v0/z1/z4/z1/z2/_1_  (.A(\v0/z1/z4/z1/temp [3]),
    .B(\v0/z1/z4/z1/temp [2]),
    .X(\v0/z1/z4/q0 [2]));
 sky130_fd_sc_hd__and2_0 \v0/z1/z4/z2/_0_  (.A(abs_b[4]),
    .B(abs_a[6]),
    .X(\v0/z1/z4/q1 [0]));
 sky130_fd_sc_hd__and2_0 \v0/z1/z4/z2/_1_  (.A(abs_b[4]),
    .B(abs_a[7]),
    .X(\v0/z1/z4/z2/temp [0]));
 sky130_fd_sc_hd__and2_0 \v0/z1/z4/z2/_2_  (.A(abs_a[6]),
    .B(abs_b[5]),
    .X(\v0/z1/z4/z2/temp [1]));
 sky130_fd_sc_hd__and2_0 \v0/z1/z4/z2/_3_  (.A(abs_a[7]),
    .B(abs_b[5]),
    .X(\v0/z1/z4/z2/temp [2]));
 sky130_fd_sc_hd__and2_0 \v0/z1/z4/z2/z1/_0_  (.A(\v0/z1/z4/z2/temp [1]),
    .B(\v0/z1/z4/z2/temp [0]),
    .X(\v0/z1/z4/z2/temp [3]));
 sky130_fd_sc_hd__xor2_1 \v0/z1/z4/z2/z1/_1_  (.A(\v0/z1/z4/z2/temp [1]),
    .B(\v0/z1/z4/z2/temp [0]),
    .X(\v0/z1/z4/q1 [1]));
 sky130_fd_sc_hd__and2_0 \v0/z1/z4/z2/z2/_0_  (.A(\v0/z1/z4/z2/temp [3]),
    .B(\v0/z1/z4/z2/temp [2]),
    .X(\v0/z1/z4/q1 [3]));
 sky130_fd_sc_hd__xor2_1 \v0/z1/z4/z2/z2/_1_  (.A(\v0/z1/z4/z2/temp [3]),
    .B(\v0/z1/z4/z2/temp [2]),
    .X(\v0/z1/z4/q1 [2]));
 sky130_fd_sc_hd__and2_0 \v0/z1/z4/z3/_0_  (.A(abs_b[6]),
    .B(abs_a[4]),
    .X(\v0/z1/z4/q2 [0]));
 sky130_fd_sc_hd__and2_0 \v0/z1/z4/z3/_1_  (.A(abs_b[6]),
    .B(abs_a[5]),
    .X(\v0/z1/z4/z3/temp [0]));
 sky130_fd_sc_hd__and2_0 \v0/z1/z4/z3/_2_  (.A(abs_a[4]),
    .B(abs_b[7]),
    .X(\v0/z1/z4/z3/temp [1]));
 sky130_fd_sc_hd__and2_0 \v0/z1/z4/z3/_3_  (.A(abs_a[5]),
    .B(abs_b[7]),
    .X(\v0/z1/z4/z3/temp [2]));
 sky130_fd_sc_hd__and2_0 \v0/z1/z4/z3/z1/_0_  (.A(\v0/z1/z4/z3/temp [1]),
    .B(\v0/z1/z4/z3/temp [0]),
    .X(\v0/z1/z4/z3/temp [3]));
 sky130_fd_sc_hd__xor2_1 \v0/z1/z4/z3/z1/_1_  (.A(\v0/z1/z4/z3/temp [1]),
    .B(\v0/z1/z4/z3/temp [0]),
    .X(\v0/z1/z4/q2 [1]));
 sky130_fd_sc_hd__and2_0 \v0/z1/z4/z3/z2/_0_  (.A(\v0/z1/z4/z3/temp [3]),
    .B(\v0/z1/z4/z3/temp [2]),
    .X(\v0/z1/z4/q2 [3]));
 sky130_fd_sc_hd__xor2_1 \v0/z1/z4/z3/z2/_1_  (.A(\v0/z1/z4/z3/temp [3]),
    .B(\v0/z1/z4/z3/temp [2]),
    .X(\v0/z1/z4/q2 [2]));
 sky130_fd_sc_hd__and2_0 \v0/z1/z4/z4/_0_  (.A(abs_b[6]),
    .B(abs_a[6]),
    .X(\v0/z1/z4/q3 [0]));
 sky130_fd_sc_hd__and2_0 \v0/z1/z4/z4/_1_  (.A(abs_b[6]),
    .B(abs_a[7]),
    .X(\v0/z1/z4/z4/temp [0]));
 sky130_fd_sc_hd__and2_0 \v0/z1/z4/z4/_2_  (.A(abs_a[6]),
    .B(abs_b[7]),
    .X(\v0/z1/z4/z4/temp [1]));
 sky130_fd_sc_hd__and2_0 \v0/z1/z4/z4/_3_  (.A(abs_a[7]),
    .B(abs_b[7]),
    .X(\v0/z1/z4/z4/temp [2]));
 sky130_fd_sc_hd__and2_0 \v0/z1/z4/z4/z1/_0_  (.A(\v0/z1/z4/z4/temp [1]),
    .B(\v0/z1/z4/z4/temp [0]),
    .X(\v0/z1/z4/z4/temp [3]));
 sky130_fd_sc_hd__xor2_1 \v0/z1/z4/z4/z1/_1_  (.A(\v0/z1/z4/z4/temp [1]),
    .B(\v0/z1/z4/z4/temp [0]),
    .X(\v0/z1/z4/q3 [1]));
 sky130_fd_sc_hd__and2_0 \v0/z1/z4/z4/z2/_0_  (.A(\v0/z1/z4/z4/temp [3]),
    .B(\v0/z1/z4/z4/temp [2]),
    .X(\v0/z1/z4/q3 [3]));
 sky130_fd_sc_hd__xor2_1 \v0/z1/z4/z4/z2/_1_  (.A(\v0/z1/z4/z4/temp [3]),
    .B(\v0/z1/z4/z4/temp [2]),
    .X(\v0/z1/z4/q3 [2]));
 sky130_fd_sc_hd__xnor2_1 \v0/z1/z4/z5/_07_  (.A(\v0/z1/z4/q0 [2]),
    .B(\v0/z1/z4/q1 [0]),
    .Y(\v0/z1/z4/z5/_00_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z1/z4/z5/_08_  (.A(\v0/z1/z4/_02_ ),
    .B(\v0/z1/z4/z5/_00_ ),
    .Y(\v0/z1/z4/q4 [0]));
 sky130_fd_sc_hd__maj3_1 \v0/z1/z4/z5/_09_  (.A(\v0/z1/z4/q0 [2]),
    .B(\v0/z1/z4/q1 [0]),
    .C(\v0/z1/z4/_02_ ),
    .X(\v0/z1/z4/z5/_01_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z1/z4/z5/_10_  (.A(\v0/z1/z4/q0 [3]),
    .B(\v0/z1/z4/q1 [1]),
    .Y(\v0/z1/z4/z5/_02_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z1/z4/z5/_11_  (.A(\v0/z1/z4/z5/_01_ ),
    .B(\v0/z1/z4/z5/_02_ ),
    .Y(\v0/z1/z4/q4 [1]));
 sky130_fd_sc_hd__maj3_1 \v0/z1/z4/z5/_12_  (.A(\v0/z1/z4/q0 [3]),
    .B(\v0/z1/z4/q1 [1]),
    .C(\v0/z1/z4/z5/_01_ ),
    .X(\v0/z1/z4/z5/_03_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z1/z4/z5/_13_  (.A(\v0/z1/z4/_00_ ),
    .B(\v0/z1/z4/q1 [2]),
    .Y(\v0/z1/z4/z5/_04_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z1/z4/z5/_14_  (.A(\v0/z1/z4/z5/_03_ ),
    .B(\v0/z1/z4/z5/_04_ ),
    .Y(\v0/z1/z4/q4 [2]));
 sky130_fd_sc_hd__maj3_1 \v0/z1/z4/z5/_15_  (.A(\v0/z1/z4/_00_ ),
    .B(\v0/z1/z4/q1 [2]),
    .C(\v0/z1/z4/z5/_03_ ),
    .X(\v0/z1/z4/z5/_05_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z1/z4/z5/_16_  (.A(\v0/z1/z4/_01_ ),
    .B(\v0/z1/z4/q1 [3]),
    .Y(\v0/z1/z4/z5/_06_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z1/z4/z5/_17_  (.A(\v0/z1/z4/z5/_05_ ),
    .B(\v0/z1/z4/z5/_06_ ),
    .Y(\v0/z1/z4/q4 [3]));
 sky130_fd_sc_hd__maj3_1 \v0/z1/z4/z5/_18_  (.A(\v0/z1/z4/_01_ ),
    .B(\v0/z1/z4/q1 [3]),
    .C(\v0/z1/z4/z5/_05_ ),
    .X(\v0/z1/z4/z5/Cout ));
 sky130_fd_sc_hd__xnor2_1 \v0/z1/z4/z6/_19_  (.A(\v0/z1/z4/_05_ ),
    .B(\v0/z1/z4/q2 [0]),
    .Y(\v0/z1/z4/z6/_00_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z1/z4/z6/_20_  (.A(\v0/z1/z4/_07_ ),
    .B(\v0/z1/z4/z6/_00_ ),
    .Y(\v0/z1/z4/q5 [0]));
 sky130_fd_sc_hd__maj3_1 \v0/z1/z4/z6/_21_  (.A(\v0/z1/z4/_05_ ),
    .B(\v0/z1/z4/q2 [0]),
    .C(\v0/z1/z4/_07_ ),
    .X(\v0/z1/z4/z6/_01_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z1/z4/z6/_22_  (.A(\v0/z1/z4/_06_ ),
    .B(\v0/z1/z4/q2 [1]),
    .Y(\v0/z1/z4/z6/_02_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z1/z4/z6/_23_  (.A(\v0/z1/z4/z6/_01_ ),
    .B(\v0/z1/z4/z6/_02_ ),
    .Y(\v0/z1/z4/q5 [1]));
 sky130_fd_sc_hd__maj3_1 \v0/z1/z4/z6/_24_  (.A(\v0/z1/z4/_06_ ),
    .B(\v0/z1/z4/q2 [1]),
    .C(\v0/z1/z4/z6/_01_ ),
    .X(\v0/z1/z4/z6/_03_ ));
 sky130_fd_sc_hd__lpflow_inputiso1p_1 \v0/z1/z4/z6/_25_  (.A(\v0/z1/z4/q3 [0]),
    .SLEEP(\v0/z1/z4/q2 [2]),
    .X(\v0/z1/z4/z6/_04_ ));
 sky130_fd_sc_hd__and2_0 \v0/z1/z4/z6/_26_  (.A(\v0/z1/z4/q3 [0]),
    .B(\v0/z1/z4/q2 [2]),
    .X(\v0/z1/z4/z6/_05_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z1/z4/z6/_27_  (.A(\v0/z1/z4/q3 [0]),
    .B(\v0/z1/z4/q2 [2]),
    .Y(\v0/z1/z4/z6/_06_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z1/z4/z6/_28_  (.A(\v0/z1/z4/z6/_04_ ),
    .B(\v0/z1/z4/z6/_06_ ),
    .Y(\v0/z1/z4/z6/_07_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z1/z4/z6/_29_  (.A(\v0/z1/z4/z6/_03_ ),
    .B(\v0/z1/z4/z6/_07_ ),
    .Y(\v0/z1/z4/q5 [2]));
 sky130_fd_sc_hd__nand2_1 \v0/z1/z4/z6/_30_  (.A(\v0/z1/z4/q3 [1]),
    .B(\v0/z1/z4/q2 [3]),
    .Y(\v0/z1/z4/z6/_08_ ));
 sky130_fd_sc_hd__xor2_1 \v0/z1/z4/z6/_31_  (.A(\v0/z1/z4/q3 [1]),
    .B(\v0/z1/z4/q2 [3]),
    .X(\v0/z1/z4/z6/_09_ ));
 sky130_fd_sc_hd__o21ai_0 \v0/z1/z4/z6/_32_  (.A1(\v0/z1/z4/z6/_03_ ),
    .A2(\v0/z1/z4/z6/_05_ ),
    .B1(\v0/z1/z4/z6/_04_ ),
    .Y(\v0/z1/z4/z6/_10_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z1/z4/z6/_33_  (.A(\v0/z1/z4/z6/_09_ ),
    .B(\v0/z1/z4/z6/_10_ ),
    .Y(\v0/z1/z4/q5 [3]));
 sky130_fd_sc_hd__nor2_1 \v0/z1/z4/z6/_34_  (.A(\v0/z1/z4/q3 [2]),
    .B(\v0/z1/z4/_03_ ),
    .Y(\v0/z1/z4/z6/_11_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z1/z4/z6/_35_  (.A(\v0/z1/z4/q3 [2]),
    .B(\v0/z1/z4/_03_ ),
    .Y(\v0/z1/z4/z6/_12_ ));
 sky130_fd_sc_hd__nand2b_1 \v0/z1/z4/z6/_36_  (.A_N(\v0/z1/z4/z6/_11_ ),
    .B(\v0/z1/z4/z6/_12_ ),
    .Y(\v0/z1/z4/z6/_13_ ));
 sky130_fd_sc_hd__o221ai_1 \v0/z1/z4/z6/_37_  (.A1(\v0/z1/z4/q3 [1]),
    .A2(\v0/z1/z4/q2 [3]),
    .B1(\v0/z1/z4/z6/_03_ ),
    .B2(\v0/z1/z4/z6/_05_ ),
    .C1(\v0/z1/z4/z6/_04_ ),
    .Y(\v0/z1/z4/z6/_14_ ));
 sky130_fd_sc_hd__a21oi_1 \v0/z1/z4/z6/_38_  (.A1(\v0/z1/z4/z6/_08_ ),
    .A2(\v0/z1/z4/z6/_14_ ),
    .B1(\v0/z1/z4/z6/_13_ ),
    .Y(\v0/z1/z4/z6/_15_ ));
 sky130_fd_sc_hd__and3_1 \v0/z1/z4/z6/_39_  (.A(\v0/z1/z4/z6/_08_ ),
    .B(\v0/z1/z4/z6/_13_ ),
    .C(\v0/z1/z4/z6/_14_ ),
    .X(\v0/z1/z4/z6/_16_ ));
 sky130_fd_sc_hd__nor2_1 \v0/z1/z4/z6/_40_  (.A(\v0/z1/z4/z6/_15_ ),
    .B(\v0/z1/z4/z6/_16_ ),
    .Y(\v0/z1/z4/q5 [4]));
 sky130_fd_sc_hd__xnor2_1 \v0/z1/z4/z6/_41_  (.A(\v0/z1/z4/q3 [3]),
    .B(\v0/z1/z4/_04_ ),
    .Y(\v0/z1/z4/z6/_17_ ));
 sky130_fd_sc_hd__a31oi_1 \v0/z1/z4/z6/_42_  (.A1(\v0/z1/z4/z6/_08_ ),
    .A2(\v0/z1/z4/z6/_12_ ),
    .A3(\v0/z1/z4/z6/_14_ ),
    .B1(\v0/z1/z4/z6/_11_ ),
    .Y(\v0/z1/z4/z6/_18_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z1/z4/z6/_43_  (.A(\v0/z1/z4/z6/_17_ ),
    .B(\v0/z1/z4/z6/_18_ ),
    .Y(\v0/z1/z4/q5 [5]));
 sky130_fd_sc_hd__maj3_1 \v0/z1/z4/z6/_44_  (.A(\v0/z1/z4/q3 [3]),
    .B(\v0/z1/z4/_04_ ),
    .C(\v0/z1/z4/z6/_18_ ),
    .X(\v0/z1/z4/z6/Cout ));
 sky130_fd_sc_hd__xnor2_1 \v0/z1/z4/z7/_19_  (.A(\v0/z1/z4/q5 [0]),
    .B(\v0/z1/z4/q4 [0]),
    .Y(\v0/z1/z4/z7/_00_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z1/z4/z7/_20_  (.A(\v0/z1/z4/_10_ ),
    .B(\v0/z1/z4/z7/_00_ ),
    .Y(\v0/z1/q3 [2]));
 sky130_fd_sc_hd__maj3_1 \v0/z1/z4/z7/_21_  (.A(\v0/z1/z4/q5 [0]),
    .B(\v0/z1/z4/q4 [0]),
    .C(\v0/z1/z4/_10_ ),
    .X(\v0/z1/z4/z7/_01_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z1/z4/z7/_22_  (.A(\v0/z1/z4/q5 [1]),
    .B(\v0/z1/z4/q4 [1]),
    .Y(\v0/z1/z4/z7/_02_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z1/z4/z7/_23_  (.A(\v0/z1/z4/z7/_01_ ),
    .B(\v0/z1/z4/z7/_02_ ),
    .Y(\v0/z1/q3 [3]));
 sky130_fd_sc_hd__maj3_1 \v0/z1/z4/z7/_24_  (.A(\v0/z1/z4/q5 [1]),
    .B(\v0/z1/z4/q4 [1]),
    .C(\v0/z1/z4/z7/_01_ ),
    .X(\v0/z1/z4/z7/_03_ ));
 sky130_fd_sc_hd__lpflow_inputiso1p_1 \v0/z1/z4/z7/_25_  (.A(\v0/z1/z4/q5 [2]),
    .SLEEP(\v0/z1/z4/q4 [2]),
    .X(\v0/z1/z4/z7/_04_ ));
 sky130_fd_sc_hd__and2_0 \v0/z1/z4/z7/_26_  (.A(\v0/z1/z4/q5 [2]),
    .B(\v0/z1/z4/q4 [2]),
    .X(\v0/z1/z4/z7/_05_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z1/z4/z7/_27_  (.A(\v0/z1/z4/q5 [2]),
    .B(\v0/z1/z4/q4 [2]),
    .Y(\v0/z1/z4/z7/_06_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z1/z4/z7/_28_  (.A(\v0/z1/z4/z7/_04_ ),
    .B(\v0/z1/z4/z7/_06_ ),
    .Y(\v0/z1/z4/z7/_07_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z1/z4/z7/_29_  (.A(\v0/z1/z4/z7/_03_ ),
    .B(\v0/z1/z4/z7/_07_ ),
    .Y(\v0/z1/q3 [4]));
 sky130_fd_sc_hd__nand2_1 \v0/z1/z4/z7/_30_  (.A(\v0/z1/z4/q5 [3]),
    .B(\v0/z1/z4/q4 [3]),
    .Y(\v0/z1/z4/z7/_08_ ));
 sky130_fd_sc_hd__xor2_1 \v0/z1/z4/z7/_31_  (.A(\v0/z1/z4/q5 [3]),
    .B(\v0/z1/z4/q4 [3]),
    .X(\v0/z1/z4/z7/_09_ ));
 sky130_fd_sc_hd__o21ai_0 \v0/z1/z4/z7/_32_  (.A1(\v0/z1/z4/z7/_03_ ),
    .A2(\v0/z1/z4/z7/_05_ ),
    .B1(\v0/z1/z4/z7/_04_ ),
    .Y(\v0/z1/z4/z7/_10_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z1/z4/z7/_33_  (.A(\v0/z1/z4/z7/_09_ ),
    .B(\v0/z1/z4/z7/_10_ ),
    .Y(\v0/z1/q3 [5]));
 sky130_fd_sc_hd__nor2_1 \v0/z1/z4/z7/_34_  (.A(\v0/z1/z4/q5 [4]),
    .B(\v0/z1/z4/_08_ ),
    .Y(\v0/z1/z4/z7/_11_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z1/z4/z7/_35_  (.A(\v0/z1/z4/q5 [4]),
    .B(\v0/z1/z4/_08_ ),
    .Y(\v0/z1/z4/z7/_12_ ));
 sky130_fd_sc_hd__nand2b_1 \v0/z1/z4/z7/_36_  (.A_N(\v0/z1/z4/z7/_11_ ),
    .B(\v0/z1/z4/z7/_12_ ),
    .Y(\v0/z1/z4/z7/_13_ ));
 sky130_fd_sc_hd__o221ai_1 \v0/z1/z4/z7/_37_  (.A1(\v0/z1/z4/q5 [3]),
    .A2(\v0/z1/z4/q4 [3]),
    .B1(\v0/z1/z4/z7/_03_ ),
    .B2(\v0/z1/z4/z7/_05_ ),
    .C1(\v0/z1/z4/z7/_04_ ),
    .Y(\v0/z1/z4/z7/_14_ ));
 sky130_fd_sc_hd__a21oi_1 \v0/z1/z4/z7/_38_  (.A1(\v0/z1/z4/z7/_08_ ),
    .A2(\v0/z1/z4/z7/_14_ ),
    .B1(\v0/z1/z4/z7/_13_ ),
    .Y(\v0/z1/z4/z7/_15_ ));
 sky130_fd_sc_hd__and3_1 \v0/z1/z4/z7/_39_  (.A(\v0/z1/z4/z7/_08_ ),
    .B(\v0/z1/z4/z7/_13_ ),
    .C(\v0/z1/z4/z7/_14_ ),
    .X(\v0/z1/z4/z7/_16_ ));
 sky130_fd_sc_hd__nor2_1 \v0/z1/z4/z7/_40_  (.A(\v0/z1/z4/z7/_15_ ),
    .B(\v0/z1/z4/z7/_16_ ),
    .Y(\v0/z1/q3 [6]));
 sky130_fd_sc_hd__xnor2_1 \v0/z1/z4/z7/_41_  (.A(\v0/z1/z4/q5 [5]),
    .B(\v0/z1/z4/_09_ ),
    .Y(\v0/z1/z4/z7/_17_ ));
 sky130_fd_sc_hd__a31oi_1 \v0/z1/z4/z7/_42_  (.A1(\v0/z1/z4/z7/_08_ ),
    .A2(\v0/z1/z4/z7/_12_ ),
    .A3(\v0/z1/z4/z7/_14_ ),
    .B1(\v0/z1/z4/z7/_11_ ),
    .Y(\v0/z1/z4/z7/_18_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z1/z4/z7/_43_  (.A(\v0/z1/z4/z7/_17_ ),
    .B(\v0/z1/z4/z7/_18_ ),
    .Y(\v0/z1/q3 [7]));
 sky130_fd_sc_hd__maj3_1 \v0/z1/z4/z7/_44_  (.A(\v0/z1/z4/q5 [5]),
    .B(\v0/z1/z4/_09_ ),
    .C(\v0/z1/z4/z7/_18_ ),
    .X(\v0/z1/z4/z7/Cout ));
 sky130_fd_sc_hd__xnor2_1 \v0/z1/z5/_27_  (.A(\v0/z1/q0 [4]),
    .B(\v0/z1/q1 [0]),
    .Y(\v0/z1/z5/_00_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z1/z5/_28_  (.A(\v0/z1/_04_ ),
    .B(\v0/z1/z5/_00_ ),
    .Y(\v0/z1/q4 [0]));
 sky130_fd_sc_hd__maj3_1 \v0/z1/z5/_29_  (.A(\v0/z1/q0 [4]),
    .B(\v0/z1/q1 [0]),
    .C(\v0/z1/_04_ ),
    .X(\v0/z1/z5/_01_ ));
 sky130_fd_sc_hd__lpflow_inputiso1p_1 \v0/z1/z5/_30_  (.A(\v0/z1/q0 [5]),
    .SLEEP(\v0/z1/q1 [1]),
    .X(\v0/z1/z5/_02_ ));
 sky130_fd_sc_hd__and2_0 \v0/z1/z5/_31_  (.A(\v0/z1/q0 [5]),
    .B(\v0/z1/q1 [1]),
    .X(\v0/z1/z5/_03_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z1/z5/_32_  (.A(\v0/z1/q0 [5]),
    .B(\v0/z1/q1 [1]),
    .Y(\v0/z1/z5/_04_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z1/z5/_33_  (.A(\v0/z1/z5/_02_ ),
    .B(\v0/z1/z5/_04_ ),
    .Y(\v0/z1/z5/_05_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z1/z5/_34_  (.A(\v0/z1/z5/_01_ ),
    .B(\v0/z1/z5/_05_ ),
    .Y(\v0/z1/q4 [1]));
 sky130_fd_sc_hd__nand2_1 \v0/z1/z5/_35_  (.A(\v0/z1/q0 [6]),
    .B(\v0/z1/q1 [2]),
    .Y(\v0/z1/z5/_06_ ));
 sky130_fd_sc_hd__xor2_1 \v0/z1/z5/_36_  (.A(\v0/z1/q0 [6]),
    .B(\v0/z1/q1 [2]),
    .X(\v0/z1/z5/_07_ ));
 sky130_fd_sc_hd__o21ai_0 \v0/z1/z5/_37_  (.A1(\v0/z1/z5/_01_ ),
    .A2(\v0/z1/z5/_03_ ),
    .B1(\v0/z1/z5/_02_ ),
    .Y(\v0/z1/z5/_08_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z1/z5/_38_  (.A(\v0/z1/z5/_07_ ),
    .B(\v0/z1/z5/_08_ ),
    .Y(\v0/z1/q4 [2]));
 sky130_fd_sc_hd__nor2_1 \v0/z1/z5/_39_  (.A(\v0/z1/q0 [7]),
    .B(\v0/z1/q1 [3]),
    .Y(\v0/z1/z5/_09_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z1/z5/_40_  (.A(\v0/z1/q0 [7]),
    .B(\v0/z1/q1 [3]),
    .Y(\v0/z1/z5/_10_ ));
 sky130_fd_sc_hd__nor2b_1 \v0/z1/z5/_41_  (.A(\v0/z1/z5/_09_ ),
    .B_N(\v0/z1/z5/_10_ ),
    .Y(\v0/z1/z5/_11_ ));
 sky130_fd_sc_hd__o221ai_1 \v0/z1/z5/_42_  (.A1(\v0/z1/q0 [6]),
    .A2(\v0/z1/q1 [2]),
    .B1(\v0/z1/z5/_01_ ),
    .B2(\v0/z1/z5/_03_ ),
    .C1(\v0/z1/z5/_02_ ),
    .Y(\v0/z1/z5/_12_ ));
 sky130_fd_sc_hd__and2_0 \v0/z1/z5/_43_  (.A(\v0/z1/z5/_06_ ),
    .B(\v0/z1/z5/_12_ ),
    .X(\v0/z1/z5/_13_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z1/z5/_44_  (.A(\v0/z1/z5/_11_ ),
    .B(\v0/z1/z5/_13_ ),
    .Y(\v0/z1/q4 [3]));
 sky130_fd_sc_hd__nor2_1 \v0/z1/z5/_45_  (.A(\v0/z1/_00_ ),
    .B(\v0/z1/q1 [4]),
    .Y(\v0/z1/z5/_14_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z1/z5/_46_  (.A(\v0/z1/_00_ ),
    .B(\v0/z1/q1 [4]),
    .Y(\v0/z1/z5/_15_ ));
 sky130_fd_sc_hd__nand2b_1 \v0/z1/z5/_47_  (.A_N(\v0/z1/z5/_14_ ),
    .B(\v0/z1/z5/_15_ ),
    .Y(\v0/z1/z5/_16_ ));
 sky130_fd_sc_hd__a21oi_1 \v0/z1/z5/_48_  (.A1(\v0/z1/z5/_10_ ),
    .A2(\v0/z1/z5/_13_ ),
    .B1(\v0/z1/z5/_09_ ),
    .Y(\v0/z1/z5/_17_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z1/z5/_49_  (.A(\v0/z1/z5/_16_ ),
    .B(\v0/z1/z5/_17_ ),
    .Y(\v0/z1/q4 [4]));
 sky130_fd_sc_hd__a311o_1 \v0/z1/z5/_50_  (.A1(\v0/z1/z5/_06_ ),
    .A2(\v0/z1/z5/_10_ ),
    .A3(\v0/z1/z5/_12_ ),
    .B1(\v0/z1/z5/_14_ ),
    .C1(\v0/z1/z5/_09_ ),
    .X(\v0/z1/z5/_18_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z1/z5/_51_  (.A(\v0/z1/z5/_15_ ),
    .B(\v0/z1/z5/_18_ ),
    .Y(\v0/z1/z5/_19_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z1/z5/_52_  (.A(\v0/z1/_01_ ),
    .B(\v0/z1/q1 [5]),
    .Y(\v0/z1/z5/_20_ ));
 sky130_fd_sc_hd__nor2_1 \v0/z1/z5/_53_  (.A(\v0/z1/_01_ ),
    .B(\v0/z1/q1 [5]),
    .Y(\v0/z1/z5/_21_ ));
 sky130_fd_sc_hd__a31oi_1 \v0/z1/z5/_54_  (.A1(\v0/z1/z5/_15_ ),
    .A2(\v0/z1/z5/_18_ ),
    .A3(\v0/z1/z5/_20_ ),
    .B1(\v0/z1/z5/_21_ ),
    .Y(\v0/z1/z5/_22_ ));
 sky130_fd_sc_hd__a21bo_1 \v0/z1/z5/_55_  (.A1(\v0/z1/z5/_20_ ),
    .A2(\v0/z1/z5/_22_ ),
    .B1_N(\v0/z1/z5/_19_ ),
    .X(\v0/z1/z5/_23_ ));
 sky130_fd_sc_hd__o21ai_0 \v0/z1/z5/_56_  (.A1(\v0/z1/z5/_21_ ),
    .A2(\v0/z1/z5/_22_ ),
    .B1(\v0/z1/z5/_23_ ),
    .Y(\v0/z1/q4 [5]));
 sky130_fd_sc_hd__xnor2_1 \v0/z1/z5/_57_  (.A(\v0/z1/_02_ ),
    .B(\v0/z1/q1 [6]),
    .Y(\v0/z1/z5/_24_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z1/z5/_58_  (.A(\v0/z1/z5/_22_ ),
    .B(\v0/z1/z5/_24_ ),
    .Y(\v0/z1/q4 [6]));
 sky130_fd_sc_hd__xnor2_1 \v0/z1/z5/_59_  (.A(\v0/z1/_03_ ),
    .B(\v0/z1/q1 [7]),
    .Y(\v0/z1/z5/_25_ ));
 sky130_fd_sc_hd__maj3_1 \v0/z1/z5/_60_  (.A(\v0/z1/_02_ ),
    .B(\v0/z1/q1 [6]),
    .C(\v0/z1/z5/_22_ ),
    .X(\v0/z1/z5/_26_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z1/z5/_61_  (.A(\v0/z1/z5/_25_ ),
    .B(\v0/z1/z5/_26_ ),
    .Y(\v0/z1/q4 [7]));
 sky130_fd_sc_hd__maj3_1 \v0/z1/z5/_62_  (.A(\v0/z1/_03_ ),
    .B(\v0/z1/q1 [7]),
    .C(\v0/z1/z5/_26_ ),
    .X(\v0/z1/z5/Cout ));
 sky130_fd_sc_hd__xnor2_1 \v0/z1/z6/_050_  (.A(\v0/z1/_09_ ),
    .B(\v0/z1/q2 [0]),
    .Y(\v0/z1/z6/_000_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z1/z6/_051_  (.A(\v0/z1/_13_ ),
    .B(\v0/z1/z6/_000_ ),
    .Y(\v0/z1/q5 [0]));
 sky130_fd_sc_hd__maj3_1 \v0/z1/z6/_052_  (.A(\v0/z1/_09_ ),
    .B(\v0/z1/q2 [0]),
    .C(\v0/z1/_13_ ),
    .X(\v0/z1/z6/_001_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z1/z6/_053_  (.A(\v0/z1/_10_ ),
    .B(\v0/z1/q2 [1]),
    .Y(\v0/z1/z6/_002_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z1/z6/_054_  (.A(\v0/z1/z6/_001_ ),
    .B(\v0/z1/z6/_002_ ),
    .Y(\v0/z1/q5 [1]));
 sky130_fd_sc_hd__maj3_1 \v0/z1/z6/_055_  (.A(\v0/z1/_10_ ),
    .B(\v0/z1/q2 [1]),
    .C(\v0/z1/z6/_001_ ),
    .X(\v0/z1/z6/_003_ ));
 sky130_fd_sc_hd__lpflow_inputiso1p_1 \v0/z1/z6/_056_  (.A(\v0/z1/_11_ ),
    .SLEEP(\v0/z1/q2 [2]),
    .X(\v0/z1/z6/_004_ ));
 sky130_fd_sc_hd__and2_0 \v0/z1/z6/_057_  (.A(\v0/z1/_11_ ),
    .B(\v0/z1/q2 [2]),
    .X(\v0/z1/z6/_005_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z1/z6/_058_  (.A(\v0/z1/_11_ ),
    .B(\v0/z1/q2 [2]),
    .Y(\v0/z1/z6/_006_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z1/z6/_059_  (.A(\v0/z1/z6/_004_ ),
    .B(\v0/z1/z6/_006_ ),
    .Y(\v0/z1/z6/_007_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z1/z6/_060_  (.A(\v0/z1/z6/_003_ ),
    .B(\v0/z1/z6/_007_ ),
    .Y(\v0/z1/q5 [2]));
 sky130_fd_sc_hd__nor2_1 \v0/z1/z6/_061_  (.A(\v0/z1/_12_ ),
    .B(\v0/z1/q2 [3]),
    .Y(\v0/z1/z6/_008_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z1/z6/_062_  (.A(\v0/z1/_12_ ),
    .B(\v0/z1/q2 [3]),
    .Y(\v0/z1/z6/_009_ ));
 sky130_fd_sc_hd__clkinv_1 \v0/z1/z6/_063_  (.A(\v0/z1/z6/_009_ ),
    .Y(\v0/z1/z6/_010_ ));
 sky130_fd_sc_hd__nor2_1 \v0/z1/z6/_064_  (.A(\v0/z1/z6/_008_ ),
    .B(\v0/z1/z6/_010_ ),
    .Y(\v0/z1/z6/_011_ ));
 sky130_fd_sc_hd__o21ai_0 \v0/z1/z6/_065_  (.A1(\v0/z1/z6/_003_ ),
    .A2(\v0/z1/z6/_005_ ),
    .B1(\v0/z1/z6/_004_ ),
    .Y(\v0/z1/z6/_012_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z1/z6/_066_  (.A(\v0/z1/z6/_011_ ),
    .B(\v0/z1/z6/_012_ ),
    .Y(\v0/z1/q5 [3]));
 sky130_fd_sc_hd__lpflow_inputiso1p_1 \v0/z1/z6/_067_  (.A(\v0/z1/q3 [0]),
    .SLEEP(\v0/z1/q2 [4]),
    .X(\v0/z1/z6/_013_ ));
 sky130_fd_sc_hd__and2_0 \v0/z1/z6/_068_  (.A(\v0/z1/q3 [0]),
    .B(\v0/z1/q2 [4]),
    .X(\v0/z1/z6/_014_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z1/z6/_069_  (.A(\v0/z1/q3 [0]),
    .B(\v0/z1/q2 [4]),
    .Y(\v0/z1/z6/_015_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z1/z6/_070_  (.A(\v0/z1/z6/_013_ ),
    .B(\v0/z1/z6/_015_ ),
    .Y(\v0/z1/z6/_016_ ));
 sky130_fd_sc_hd__o221a_1 \v0/z1/z6/_071_  (.A1(\v0/z1/_12_ ),
    .A2(\v0/z1/q2 [3]),
    .B1(\v0/z1/z6/_003_ ),
    .B2(\v0/z1/z6/_005_ ),
    .C1(\v0/z1/z6/_004_ ),
    .X(\v0/z1/z6/_017_ ));
 sky130_fd_sc_hd__a21oi_1 \v0/z1/z6/_072_  (.A1(\v0/z1/z6/_009_ ),
    .A2(\v0/z1/z6/_012_ ),
    .B1(\v0/z1/z6/_008_ ),
    .Y(\v0/z1/z6/_018_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z1/z6/_073_  (.A(\v0/z1/z6/_016_ ),
    .B(\v0/z1/z6/_018_ ),
    .Y(\v0/z1/q5 [4]));
 sky130_fd_sc_hd__lpflow_inputiso1p_1 \v0/z1/z6/_074_  (.A(\v0/z1/q3 [1]),
    .SLEEP(\v0/z1/q2 [5]),
    .X(\v0/z1/z6/_019_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z1/z6/_075_  (.A(\v0/z1/q3 [1]),
    .B(\v0/z1/q2 [5]),
    .Y(\v0/z1/z6/_020_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z1/z6/_076_  (.A(\v0/z1/z6/_019_ ),
    .B(\v0/z1/z6/_020_ ),
    .Y(\v0/z1/z6/_021_ ));
 sky130_fd_sc_hd__o21ai_0 \v0/z1/z6/_077_  (.A1(\v0/z1/z6/_014_ ),
    .A2(\v0/z1/z6/_018_ ),
    .B1(\v0/z1/z6/_013_ ),
    .Y(\v0/z1/z6/_022_ ));
 sky130_fd_sc_hd__xor2_1 \v0/z1/z6/_078_  (.A(\v0/z1/z6/_021_ ),
    .B(\v0/z1/z6/_022_ ),
    .X(\v0/z1/q5 [5]));
 sky130_fd_sc_hd__nor2_1 \v0/z1/z6/_079_  (.A(\v0/z1/q3 [2]),
    .B(\v0/z1/q2 [6]),
    .Y(\v0/z1/z6/_023_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z1/z6/_080_  (.A(\v0/z1/q3 [2]),
    .B(\v0/z1/q2 [6]),
    .Y(\v0/z1/z6/_024_ ));
 sky130_fd_sc_hd__nor2b_1 \v0/z1/z6/_081_  (.A(\v0/z1/z6/_023_ ),
    .B_N(\v0/z1/z6/_024_ ),
    .Y(\v0/z1/z6/_025_ ));
 sky130_fd_sc_hd__o311ai_0 \v0/z1/z6/_082_  (.A1(\v0/z1/z6/_010_ ),
    .A2(\v0/z1/z6/_014_ ),
    .A3(\v0/z1/z6/_017_ ),
    .B1(\v0/z1/z6/_019_ ),
    .C1(\v0/z1/z6/_013_ ),
    .Y(\v0/z1/z6/_026_ ));
 sky130_fd_sc_hd__and2_0 \v0/z1/z6/_083_  (.A(\v0/z1/z6/_020_ ),
    .B(\v0/z1/z6/_026_ ),
    .X(\v0/z1/z6/_027_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z1/z6/_084_  (.A(\v0/z1/z6/_025_ ),
    .B(\v0/z1/z6/_027_ ),
    .Y(\v0/z1/q5 [6]));
 sky130_fd_sc_hd__nor2_1 \v0/z1/z6/_085_  (.A(\v0/z1/q3 [3]),
    .B(\v0/z1/q2 [7]),
    .Y(\v0/z1/z6/_028_ ));
 sky130_fd_sc_hd__and2_0 \v0/z1/z6/_086_  (.A(\v0/z1/q3 [3]),
    .B(\v0/z1/q2 [7]),
    .X(\v0/z1/z6/_029_ ));
 sky130_fd_sc_hd__nor2_1 \v0/z1/z6/_087_  (.A(\v0/z1/z6/_028_ ),
    .B(\v0/z1/z6/_029_ ),
    .Y(\v0/z1/z6/_030_ ));
 sky130_fd_sc_hd__a21oi_1 \v0/z1/z6/_088_  (.A1(\v0/z1/z6/_024_ ),
    .A2(\v0/z1/z6/_027_ ),
    .B1(\v0/z1/z6/_023_ ),
    .Y(\v0/z1/z6/_031_ ));
 sky130_fd_sc_hd__xor2_1 \v0/z1/z6/_089_  (.A(\v0/z1/z6/_030_ ),
    .B(\v0/z1/z6/_031_ ),
    .X(\v0/z1/q5 [7]));
 sky130_fd_sc_hd__lpflow_inputiso1p_1 \v0/z1/z6/_090_  (.A(\v0/z1/q3 [4]),
    .SLEEP(\v0/z1/_05_ ),
    .X(\v0/z1/z6/_032_ ));
 sky130_fd_sc_hd__and2_0 \v0/z1/z6/_091_  (.A(\v0/z1/q3 [4]),
    .B(\v0/z1/_05_ ),
    .X(\v0/z1/z6/_033_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z1/z6/_092_  (.A(\v0/z1/q3 [4]),
    .B(\v0/z1/_05_ ),
    .Y(\v0/z1/z6/_034_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z1/z6/_093_  (.A(\v0/z1/z6/_032_ ),
    .B(\v0/z1/z6/_034_ ),
    .Y(\v0/z1/z6/_035_ ));
 sky130_fd_sc_hd__a311oi_1 \v0/z1/z6/_094_  (.A1(\v0/z1/z6/_020_ ),
    .A2(\v0/z1/z6/_024_ ),
    .A3(\v0/z1/z6/_026_ ),
    .B1(\v0/z1/z6/_028_ ),
    .C1(\v0/z1/z6/_023_ ),
    .Y(\v0/z1/z6/_036_ ));
 sky130_fd_sc_hd__lpflow_inputiso1p_1 \v0/z1/z6/_095_  (.A(\v0/z1/z6/_029_ ),
    .SLEEP(\v0/z1/z6/_036_ ),
    .X(\v0/z1/z6/_037_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z1/z6/_096_  (.A(\v0/z1/z6/_035_ ),
    .B(\v0/z1/z6/_037_ ),
    .Y(\v0/z1/q5 [8]));
 sky130_fd_sc_hd__lpflow_inputiso1p_1 \v0/z1/z6/_097_  (.A(\v0/z1/q3 [5]),
    .SLEEP(\v0/z1/_06_ ),
    .X(\v0/z1/z6/_038_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z1/z6/_098_  (.A(\v0/z1/q3 [5]),
    .B(\v0/z1/_06_ ),
    .Y(\v0/z1/z6/_039_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z1/z6/_099_  (.A(\v0/z1/z6/_038_ ),
    .B(\v0/z1/z6/_039_ ),
    .Y(\v0/z1/z6/_040_ ));
 sky130_fd_sc_hd__o21ai_0 \v0/z1/z6/_100_  (.A1(\v0/z1/z6/_033_ ),
    .A2(\v0/z1/z6/_037_ ),
    .B1(\v0/z1/z6/_032_ ),
    .Y(\v0/z1/z6/_041_ ));
 sky130_fd_sc_hd__xor2_1 \v0/z1/z6/_101_  (.A(\v0/z1/z6/_040_ ),
    .B(\v0/z1/z6/_041_ ),
    .X(\v0/z1/q5 [9]));
 sky130_fd_sc_hd__nor2_1 \v0/z1/z6/_102_  (.A(\v0/z1/q3 [6]),
    .B(\v0/z1/_07_ ),
    .Y(\v0/z1/z6/_042_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z1/z6/_103_  (.A(\v0/z1/q3 [6]),
    .B(\v0/z1/_07_ ),
    .Y(\v0/z1/z6/_043_ ));
 sky130_fd_sc_hd__nand2b_1 \v0/z1/z6/_104_  (.A_N(\v0/z1/z6/_042_ ),
    .B(\v0/z1/z6/_043_ ),
    .Y(\v0/z1/z6/_044_ ));
 sky130_fd_sc_hd__o311ai_0 \v0/z1/z6/_105_  (.A1(\v0/z1/z6/_029_ ),
    .A2(\v0/z1/z6/_033_ ),
    .A3(\v0/z1/z6/_036_ ),
    .B1(\v0/z1/z6/_038_ ),
    .C1(\v0/z1/z6/_032_ ),
    .Y(\v0/z1/z6/_045_ ));
 sky130_fd_sc_hd__a21oi_1 \v0/z1/z6/_106_  (.A1(\v0/z1/z6/_039_ ),
    .A2(\v0/z1/z6/_045_ ),
    .B1(\v0/z1/z6/_044_ ),
    .Y(\v0/z1/z6/_046_ ));
 sky130_fd_sc_hd__and3_1 \v0/z1/z6/_107_  (.A(\v0/z1/z6/_039_ ),
    .B(\v0/z1/z6/_044_ ),
    .C(\v0/z1/z6/_045_ ),
    .X(\v0/z1/z6/_047_ ));
 sky130_fd_sc_hd__nor2_1 \v0/z1/z6/_108_  (.A(\v0/z1/z6/_046_ ),
    .B(\v0/z1/z6/_047_ ),
    .Y(\v0/z1/q5 [10]));
 sky130_fd_sc_hd__xnor2_1 \v0/z1/z6/_109_  (.A(\v0/z1/q3 [7]),
    .B(\v0/z1/_08_ ),
    .Y(\v0/z1/z6/_048_ ));
 sky130_fd_sc_hd__a31oi_1 \v0/z1/z6/_110_  (.A1(\v0/z1/z6/_039_ ),
    .A2(\v0/z1/z6/_043_ ),
    .A3(\v0/z1/z6/_045_ ),
    .B1(\v0/z1/z6/_042_ ),
    .Y(\v0/z1/z6/_049_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z1/z6/_111_  (.A(\v0/z1/z6/_048_ ),
    .B(\v0/z1/z6/_049_ ),
    .Y(\v0/z1/q5 [11]));
 sky130_fd_sc_hd__maj3_1 \v0/z1/z6/_112_  (.A(\v0/z1/q3 [7]),
    .B(\v0/z1/_08_ ),
    .C(\v0/z1/z6/_049_ ),
    .X(\v0/z1/z6/Cout ));
 sky130_fd_sc_hd__xnor2_1 \v0/z1/z7/_050_  (.A(\v0/z1/q5 [0]),
    .B(\v0/z1/q4 [0]),
    .Y(\v0/z1/z7/_000_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z1/z7/_051_  (.A(\v0/z1/_18_ ),
    .B(\v0/z1/z7/_000_ ),
    .Y(unsign[4]));
 sky130_fd_sc_hd__maj3_1 \v0/z1/z7/_052_  (.A(\v0/z1/q5 [0]),
    .B(\v0/z1/q4 [0]),
    .C(\v0/z1/_18_ ),
    .X(\v0/z1/z7/_001_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z1/z7/_053_  (.A(\v0/z1/q5 [1]),
    .B(\v0/z1/q4 [1]),
    .Y(\v0/z1/z7/_002_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z1/z7/_054_  (.A(\v0/z1/z7/_001_ ),
    .B(\v0/z1/z7/_002_ ),
    .Y(unsign[5]));
 sky130_fd_sc_hd__maj3_1 \v0/z1/z7/_055_  (.A(\v0/z1/q5 [1]),
    .B(\v0/z1/q4 [1]),
    .C(\v0/z1/z7/_001_ ),
    .X(\v0/z1/z7/_003_ ));
 sky130_fd_sc_hd__lpflow_inputiso1p_1 \v0/z1/z7/_056_  (.A(\v0/z1/q5 [2]),
    .SLEEP(\v0/z1/q4 [2]),
    .X(\v0/z1/z7/_004_ ));
 sky130_fd_sc_hd__and2_0 \v0/z1/z7/_057_  (.A(\v0/z1/q5 [2]),
    .B(\v0/z1/q4 [2]),
    .X(\v0/z1/z7/_005_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z1/z7/_058_  (.A(\v0/z1/q5 [2]),
    .B(\v0/z1/q4 [2]),
    .Y(\v0/z1/z7/_006_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z1/z7/_059_  (.A(\v0/z1/z7/_004_ ),
    .B(\v0/z1/z7/_006_ ),
    .Y(\v0/z1/z7/_007_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z1/z7/_060_  (.A(\v0/z1/z7/_003_ ),
    .B(\v0/z1/z7/_007_ ),
    .Y(unsign[6]));
 sky130_fd_sc_hd__nor2_1 \v0/z1/z7/_061_  (.A(\v0/z1/q5 [3]),
    .B(\v0/z1/q4 [3]),
    .Y(\v0/z1/z7/_008_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z1/z7/_062_  (.A(\v0/z1/q5 [3]),
    .B(\v0/z1/q4 [3]),
    .Y(\v0/z1/z7/_009_ ));
 sky130_fd_sc_hd__clkinv_1 \v0/z1/z7/_063_  (.A(\v0/z1/z7/_009_ ),
    .Y(\v0/z1/z7/_010_ ));
 sky130_fd_sc_hd__nor2_1 \v0/z1/z7/_064_  (.A(\v0/z1/z7/_008_ ),
    .B(\v0/z1/z7/_010_ ),
    .Y(\v0/z1/z7/_011_ ));
 sky130_fd_sc_hd__o21ai_0 \v0/z1/z7/_065_  (.A1(\v0/z1/z7/_003_ ),
    .A2(\v0/z1/z7/_005_ ),
    .B1(\v0/z1/z7/_004_ ),
    .Y(\v0/z1/z7/_012_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z1/z7/_066_  (.A(\v0/z1/z7/_011_ ),
    .B(\v0/z1/z7/_012_ ),
    .Y(unsign[7]));
 sky130_fd_sc_hd__lpflow_inputiso1p_1 \v0/z1/z7/_067_  (.A(\v0/z1/q5 [4]),
    .SLEEP(\v0/z1/q4 [4]),
    .X(\v0/z1/z7/_013_ ));
 sky130_fd_sc_hd__and2_0 \v0/z1/z7/_068_  (.A(\v0/z1/q5 [4]),
    .B(\v0/z1/q4 [4]),
    .X(\v0/z1/z7/_014_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z1/z7/_069_  (.A(\v0/z1/q5 [4]),
    .B(\v0/z1/q4 [4]),
    .Y(\v0/z1/z7/_015_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z1/z7/_070_  (.A(\v0/z1/z7/_013_ ),
    .B(\v0/z1/z7/_015_ ),
    .Y(\v0/z1/z7/_016_ ));
 sky130_fd_sc_hd__o221a_1 \v0/z1/z7/_071_  (.A1(\v0/z1/q5 [3]),
    .A2(\v0/z1/q4 [3]),
    .B1(\v0/z1/z7/_003_ ),
    .B2(\v0/z1/z7/_005_ ),
    .C1(\v0/z1/z7/_004_ ),
    .X(\v0/z1/z7/_017_ ));
 sky130_fd_sc_hd__a21oi_1 \v0/z1/z7/_072_  (.A1(\v0/z1/z7/_009_ ),
    .A2(\v0/z1/z7/_012_ ),
    .B1(\v0/z1/z7/_008_ ),
    .Y(\v0/z1/z7/_018_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z1/z7/_073_  (.A(\v0/z1/z7/_016_ ),
    .B(\v0/z1/z7/_018_ ),
    .Y(\v0/q0 [8]));
 sky130_fd_sc_hd__lpflow_inputiso1p_1 \v0/z1/z7/_074_  (.A(\v0/z1/q5 [5]),
    .SLEEP(\v0/z1/q4 [5]),
    .X(\v0/z1/z7/_019_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z1/z7/_075_  (.A(\v0/z1/q5 [5]),
    .B(\v0/z1/q4 [5]),
    .Y(\v0/z1/z7/_020_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z1/z7/_076_  (.A(\v0/z1/z7/_019_ ),
    .B(\v0/z1/z7/_020_ ),
    .Y(\v0/z1/z7/_021_ ));
 sky130_fd_sc_hd__o21ai_0 \v0/z1/z7/_077_  (.A1(\v0/z1/z7/_014_ ),
    .A2(\v0/z1/z7/_018_ ),
    .B1(\v0/z1/z7/_013_ ),
    .Y(\v0/z1/z7/_022_ ));
 sky130_fd_sc_hd__xor2_1 \v0/z1/z7/_078_  (.A(\v0/z1/z7/_021_ ),
    .B(\v0/z1/z7/_022_ ),
    .X(\v0/q0 [9]));
 sky130_fd_sc_hd__nor2_1 \v0/z1/z7/_079_  (.A(\v0/z1/q5 [6]),
    .B(\v0/z1/q4 [6]),
    .Y(\v0/z1/z7/_023_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z1/z7/_080_  (.A(\v0/z1/q5 [6]),
    .B(\v0/z1/q4 [6]),
    .Y(\v0/z1/z7/_024_ ));
 sky130_fd_sc_hd__nor2b_1 \v0/z1/z7/_081_  (.A(\v0/z1/z7/_023_ ),
    .B_N(\v0/z1/z7/_024_ ),
    .Y(\v0/z1/z7/_025_ ));
 sky130_fd_sc_hd__o311ai_0 \v0/z1/z7/_082_  (.A1(\v0/z1/z7/_010_ ),
    .A2(\v0/z1/z7/_014_ ),
    .A3(\v0/z1/z7/_017_ ),
    .B1(\v0/z1/z7/_019_ ),
    .C1(\v0/z1/z7/_013_ ),
    .Y(\v0/z1/z7/_026_ ));
 sky130_fd_sc_hd__and2_0 \v0/z1/z7/_083_  (.A(\v0/z1/z7/_020_ ),
    .B(\v0/z1/z7/_026_ ),
    .X(\v0/z1/z7/_027_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z1/z7/_084_  (.A(\v0/z1/z7/_025_ ),
    .B(\v0/z1/z7/_027_ ),
    .Y(\v0/q0 [10]));
 sky130_fd_sc_hd__nor2_1 \v0/z1/z7/_085_  (.A(\v0/z1/q5 [7]),
    .B(\v0/z1/q4 [7]),
    .Y(\v0/z1/z7/_028_ ));
 sky130_fd_sc_hd__and2_0 \v0/z1/z7/_086_  (.A(\v0/z1/q5 [7]),
    .B(\v0/z1/q4 [7]),
    .X(\v0/z1/z7/_029_ ));
 sky130_fd_sc_hd__nor2_1 \v0/z1/z7/_087_  (.A(\v0/z1/z7/_028_ ),
    .B(\v0/z1/z7/_029_ ),
    .Y(\v0/z1/z7/_030_ ));
 sky130_fd_sc_hd__a21oi_1 \v0/z1/z7/_088_  (.A1(\v0/z1/z7/_024_ ),
    .A2(\v0/z1/z7/_027_ ),
    .B1(\v0/z1/z7/_023_ ),
    .Y(\v0/z1/z7/_031_ ));
 sky130_fd_sc_hd__xor2_1 \v0/z1/z7/_089_  (.A(\v0/z1/z7/_030_ ),
    .B(\v0/z1/z7/_031_ ),
    .X(\v0/q0 [11]));
 sky130_fd_sc_hd__lpflow_inputiso1p_1 \v0/z1/z7/_090_  (.A(\v0/z1/q5 [8]),
    .SLEEP(\v0/z1/_14_ ),
    .X(\v0/z1/z7/_032_ ));
 sky130_fd_sc_hd__and2_0 \v0/z1/z7/_091_  (.A(\v0/z1/q5 [8]),
    .B(\v0/z1/_14_ ),
    .X(\v0/z1/z7/_033_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z1/z7/_092_  (.A(\v0/z1/q5 [8]),
    .B(\v0/z1/_14_ ),
    .Y(\v0/z1/z7/_034_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z1/z7/_093_  (.A(\v0/z1/z7/_032_ ),
    .B(\v0/z1/z7/_034_ ),
    .Y(\v0/z1/z7/_035_ ));
 sky130_fd_sc_hd__a311oi_1 \v0/z1/z7/_094_  (.A1(\v0/z1/z7/_020_ ),
    .A2(\v0/z1/z7/_024_ ),
    .A3(\v0/z1/z7/_026_ ),
    .B1(\v0/z1/z7/_028_ ),
    .C1(\v0/z1/z7/_023_ ),
    .Y(\v0/z1/z7/_036_ ));
 sky130_fd_sc_hd__lpflow_inputiso1p_1 \v0/z1/z7/_095_  (.A(\v0/z1/z7/_029_ ),
    .SLEEP(\v0/z1/z7/_036_ ),
    .X(\v0/z1/z7/_037_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z1/z7/_096_  (.A(\v0/z1/z7/_035_ ),
    .B(\v0/z1/z7/_037_ ),
    .Y(\v0/q0 [12]));
 sky130_fd_sc_hd__lpflow_inputiso1p_1 \v0/z1/z7/_097_  (.A(\v0/z1/q5 [9]),
    .SLEEP(\v0/z1/_15_ ),
    .X(\v0/z1/z7/_038_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z1/z7/_098_  (.A(\v0/z1/q5 [9]),
    .B(\v0/z1/_15_ ),
    .Y(\v0/z1/z7/_039_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z1/z7/_099_  (.A(\v0/z1/z7/_038_ ),
    .B(\v0/z1/z7/_039_ ),
    .Y(\v0/z1/z7/_040_ ));
 sky130_fd_sc_hd__o21ai_0 \v0/z1/z7/_100_  (.A1(\v0/z1/z7/_033_ ),
    .A2(\v0/z1/z7/_037_ ),
    .B1(\v0/z1/z7/_032_ ),
    .Y(\v0/z1/z7/_041_ ));
 sky130_fd_sc_hd__xor2_1 \v0/z1/z7/_101_  (.A(\v0/z1/z7/_040_ ),
    .B(\v0/z1/z7/_041_ ),
    .X(\v0/q0 [13]));
 sky130_fd_sc_hd__nor2_1 \v0/z1/z7/_102_  (.A(\v0/z1/q5 [10]),
    .B(\v0/z1/_16_ ),
    .Y(\v0/z1/z7/_042_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z1/z7/_103_  (.A(\v0/z1/q5 [10]),
    .B(\v0/z1/_16_ ),
    .Y(\v0/z1/z7/_043_ ));
 sky130_fd_sc_hd__nand2b_1 \v0/z1/z7/_104_  (.A_N(\v0/z1/z7/_042_ ),
    .B(\v0/z1/z7/_043_ ),
    .Y(\v0/z1/z7/_044_ ));
 sky130_fd_sc_hd__o311ai_0 \v0/z1/z7/_105_  (.A1(\v0/z1/z7/_029_ ),
    .A2(\v0/z1/z7/_033_ ),
    .A3(\v0/z1/z7/_036_ ),
    .B1(\v0/z1/z7/_038_ ),
    .C1(\v0/z1/z7/_032_ ),
    .Y(\v0/z1/z7/_045_ ));
 sky130_fd_sc_hd__a21oi_1 \v0/z1/z7/_106_  (.A1(\v0/z1/z7/_039_ ),
    .A2(\v0/z1/z7/_045_ ),
    .B1(\v0/z1/z7/_044_ ),
    .Y(\v0/z1/z7/_046_ ));
 sky130_fd_sc_hd__and3_1 \v0/z1/z7/_107_  (.A(\v0/z1/z7/_039_ ),
    .B(\v0/z1/z7/_044_ ),
    .C(\v0/z1/z7/_045_ ),
    .X(\v0/z1/z7/_047_ ));
 sky130_fd_sc_hd__nor2_1 \v0/z1/z7/_108_  (.A(\v0/z1/z7/_046_ ),
    .B(\v0/z1/z7/_047_ ),
    .Y(\v0/q0 [14]));
 sky130_fd_sc_hd__xnor2_1 \v0/z1/z7/_109_  (.A(\v0/z1/q5 [11]),
    .B(\v0/z1/_17_ ),
    .Y(\v0/z1/z7/_048_ ));
 sky130_fd_sc_hd__a31oi_1 \v0/z1/z7/_110_  (.A1(\v0/z1/z7/_039_ ),
    .A2(\v0/z1/z7/_043_ ),
    .A3(\v0/z1/z7/_045_ ),
    .B1(\v0/z1/z7/_042_ ),
    .Y(\v0/z1/z7/_049_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z1/z7/_111_  (.A(\v0/z1/z7/_048_ ),
    .B(\v0/z1/z7/_049_ ),
    .Y(\v0/q0 [15]));
 sky130_fd_sc_hd__maj3_1 \v0/z1/z7/_112_  (.A(\v0/z1/q5 [11]),
    .B(\v0/z1/_17_ ),
    .C(\v0/z1/z7/_049_ ),
    .X(\v0/z1/z7/Cout ));
 sky130_fd_sc_hd__conb_1 \v0/z2/_19_  (.LO(\v0/z2/_00_ ));
 sky130_fd_sc_hd__conb_1 \v0/z2/_20_  (.LO(\v0/z2/_01_ ));
 sky130_fd_sc_hd__conb_1 \v0/z2/_21_  (.LO(\v0/z2/_02_ ));
 sky130_fd_sc_hd__conb_1 \v0/z2/_22_  (.LO(\v0/z2/_03_ ));
 sky130_fd_sc_hd__conb_1 \v0/z2/_23_  (.LO(\v0/z2/_04_ ));
 sky130_fd_sc_hd__conb_1 \v0/z2/_24_  (.LO(\v0/z2/_05_ ));
 sky130_fd_sc_hd__conb_1 \v0/z2/_25_  (.LO(\v0/z2/_06_ ));
 sky130_fd_sc_hd__conb_1 \v0/z2/_26_  (.LO(\v0/z2/_07_ ));
 sky130_fd_sc_hd__conb_1 \v0/z2/_27_  (.LO(\v0/z2/_08_ ));
 sky130_fd_sc_hd__conb_1 \v0/z2/_28_  (.LO(\v0/z2/_09_ ));
 sky130_fd_sc_hd__conb_1 \v0/z2/_29_  (.LO(\v0/z2/_10_ ));
 sky130_fd_sc_hd__conb_1 \v0/z2/_30_  (.LO(\v0/z2/_11_ ));
 sky130_fd_sc_hd__conb_1 \v0/z2/_31_  (.LO(\v0/z2/_12_ ));
 sky130_fd_sc_hd__conb_1 \v0/z2/_32_  (.LO(\v0/z2/_13_ ));
 sky130_fd_sc_hd__conb_1 \v0/z2/_33_  (.LO(\v0/z2/_14_ ));
 sky130_fd_sc_hd__conb_1 \v0/z2/_34_  (.LO(\v0/z2/_15_ ));
 sky130_fd_sc_hd__conb_1 \v0/z2/_35_  (.LO(\v0/z2/_16_ ));
 sky130_fd_sc_hd__conb_1 \v0/z2/_36_  (.LO(\v0/z2/_17_ ));
 sky130_fd_sc_hd__conb_1 \v0/z2/_37_  (.LO(\v0/z2/_18_ ));
 sky130_fd_sc_hd__conb_1 \v0/z2/z1/_11_  (.LO(\v0/z2/z1/_00_ ));
 sky130_fd_sc_hd__conb_1 \v0/z2/z1/_12_  (.LO(\v0/z2/z1/_01_ ));
 sky130_fd_sc_hd__conb_1 \v0/z2/z1/_13_  (.LO(\v0/z2/z1/_02_ ));
 sky130_fd_sc_hd__conb_1 \v0/z2/z1/_14_  (.LO(\v0/z2/z1/_03_ ));
 sky130_fd_sc_hd__conb_1 \v0/z2/z1/_15_  (.LO(\v0/z2/z1/_04_ ));
 sky130_fd_sc_hd__conb_1 \v0/z2/z1/_16_  (.LO(\v0/z2/z1/_05_ ));
 sky130_fd_sc_hd__conb_1 \v0/z2/z1/_17_  (.LO(\v0/z2/z1/_06_ ));
 sky130_fd_sc_hd__conb_1 \v0/z2/z1/_18_  (.LO(\v0/z2/z1/_07_ ));
 sky130_fd_sc_hd__conb_1 \v0/z2/z1/_19_  (.LO(\v0/z2/z1/_08_ ));
 sky130_fd_sc_hd__conb_1 \v0/z2/z1/_20_  (.LO(\v0/z2/z1/_09_ ));
 sky130_fd_sc_hd__conb_1 \v0/z2/z1/_21_  (.LO(\v0/z2/z1/_10_ ));
 sky130_fd_sc_hd__and2_0 \v0/z2/z1/z1/_0_  (.A(b[0]),
    .B(abs_a[8]),
    .X(\v0/q1 [0]));
 sky130_fd_sc_hd__and2_0 \v0/z2/z1/z1/_1_  (.A(b[0]),
    .B(abs_a[9]),
    .X(\v0/z2/z1/z1/temp [0]));
 sky130_fd_sc_hd__and2_0 \v0/z2/z1/z1/_2_  (.A(abs_a[8]),
    .B(abs_b[1]),
    .X(\v0/z2/z1/z1/temp [1]));
 sky130_fd_sc_hd__and2_0 \v0/z2/z1/z1/_3_  (.A(abs_a[9]),
    .B(abs_b[1]),
    .X(\v0/z2/z1/z1/temp [2]));
 sky130_fd_sc_hd__and2_0 \v0/z2/z1/z1/z1/_0_  (.A(\v0/z2/z1/z1/temp [1]),
    .B(\v0/z2/z1/z1/temp [0]),
    .X(\v0/z2/z1/z1/temp [3]));
 sky130_fd_sc_hd__xor2_1 \v0/z2/z1/z1/z1/_1_  (.A(\v0/z2/z1/z1/temp [1]),
    .B(\v0/z2/z1/z1/temp [0]),
    .X(\v0/q1 [1]));
 sky130_fd_sc_hd__and2_0 \v0/z2/z1/z1/z2/_0_  (.A(\v0/z2/z1/z1/temp [3]),
    .B(\v0/z2/z1/z1/temp [2]),
    .X(\v0/z2/z1/q0 [3]));
 sky130_fd_sc_hd__xor2_1 \v0/z2/z1/z1/z2/_1_  (.A(\v0/z2/z1/z1/temp [3]),
    .B(\v0/z2/z1/z1/temp [2]),
    .X(\v0/z2/z1/q0 [2]));
 sky130_fd_sc_hd__and2_0 \v0/z2/z1/z2/_0_  (.A(b[0]),
    .B(abs_a[10]),
    .X(\v0/z2/z1/q1 [0]));
 sky130_fd_sc_hd__and2_0 \v0/z2/z1/z2/_1_  (.A(b[0]),
    .B(abs_a[11]),
    .X(\v0/z2/z1/z2/temp [0]));
 sky130_fd_sc_hd__and2_0 \v0/z2/z1/z2/_2_  (.A(abs_a[10]),
    .B(abs_b[1]),
    .X(\v0/z2/z1/z2/temp [1]));
 sky130_fd_sc_hd__and2_0 \v0/z2/z1/z2/_3_  (.A(abs_a[11]),
    .B(abs_b[1]),
    .X(\v0/z2/z1/z2/temp [2]));
 sky130_fd_sc_hd__and2_0 \v0/z2/z1/z2/z1/_0_  (.A(\v0/z2/z1/z2/temp [1]),
    .B(\v0/z2/z1/z2/temp [0]),
    .X(\v0/z2/z1/z2/temp [3]));
 sky130_fd_sc_hd__xor2_1 \v0/z2/z1/z2/z1/_1_  (.A(\v0/z2/z1/z2/temp [1]),
    .B(\v0/z2/z1/z2/temp [0]),
    .X(\v0/z2/z1/q1 [1]));
 sky130_fd_sc_hd__and2_0 \v0/z2/z1/z2/z2/_0_  (.A(\v0/z2/z1/z2/temp [3]),
    .B(\v0/z2/z1/z2/temp [2]),
    .X(\v0/z2/z1/q1 [3]));
 sky130_fd_sc_hd__xor2_1 \v0/z2/z1/z2/z2/_1_  (.A(\v0/z2/z1/z2/temp [3]),
    .B(\v0/z2/z1/z2/temp [2]),
    .X(\v0/z2/z1/q1 [2]));
 sky130_fd_sc_hd__and2_0 \v0/z2/z1/z3/_0_  (.A(abs_b[2]),
    .B(abs_a[8]),
    .X(\v0/z2/z1/q2 [0]));
 sky130_fd_sc_hd__and2_0 \v0/z2/z1/z3/_1_  (.A(abs_b[2]),
    .B(abs_a[9]),
    .X(\v0/z2/z1/z3/temp [0]));
 sky130_fd_sc_hd__and2_0 \v0/z2/z1/z3/_2_  (.A(abs_a[8]),
    .B(abs_b[3]),
    .X(\v0/z2/z1/z3/temp [1]));
 sky130_fd_sc_hd__and2_0 \v0/z2/z1/z3/_3_  (.A(abs_a[9]),
    .B(abs_b[3]),
    .X(\v0/z2/z1/z3/temp [2]));
 sky130_fd_sc_hd__and2_0 \v0/z2/z1/z3/z1/_0_  (.A(\v0/z2/z1/z3/temp [1]),
    .B(\v0/z2/z1/z3/temp [0]),
    .X(\v0/z2/z1/z3/temp [3]));
 sky130_fd_sc_hd__xor2_1 \v0/z2/z1/z3/z1/_1_  (.A(\v0/z2/z1/z3/temp [1]),
    .B(\v0/z2/z1/z3/temp [0]),
    .X(\v0/z2/z1/q2 [1]));
 sky130_fd_sc_hd__and2_0 \v0/z2/z1/z3/z2/_0_  (.A(\v0/z2/z1/z3/temp [3]),
    .B(\v0/z2/z1/z3/temp [2]),
    .X(\v0/z2/z1/q2 [3]));
 sky130_fd_sc_hd__xor2_1 \v0/z2/z1/z3/z2/_1_  (.A(\v0/z2/z1/z3/temp [3]),
    .B(\v0/z2/z1/z3/temp [2]),
    .X(\v0/z2/z1/q2 [2]));
 sky130_fd_sc_hd__and2_0 \v0/z2/z1/z4/_0_  (.A(abs_b[2]),
    .B(abs_a[10]),
    .X(\v0/z2/z1/q3 [0]));
 sky130_fd_sc_hd__and2_0 \v0/z2/z1/z4/_1_  (.A(abs_b[2]),
    .B(abs_a[11]),
    .X(\v0/z2/z1/z4/temp [0]));
 sky130_fd_sc_hd__and2_0 \v0/z2/z1/z4/_2_  (.A(abs_a[10]),
    .B(abs_b[3]),
    .X(\v0/z2/z1/z4/temp [1]));
 sky130_fd_sc_hd__and2_0 \v0/z2/z1/z4/_3_  (.A(abs_a[11]),
    .B(abs_b[3]),
    .X(\v0/z2/z1/z4/temp [2]));
 sky130_fd_sc_hd__and2_0 \v0/z2/z1/z4/z1/_0_  (.A(\v0/z2/z1/z4/temp [1]),
    .B(\v0/z2/z1/z4/temp [0]),
    .X(\v0/z2/z1/z4/temp [3]));
 sky130_fd_sc_hd__xor2_1 \v0/z2/z1/z4/z1/_1_  (.A(\v0/z2/z1/z4/temp [1]),
    .B(\v0/z2/z1/z4/temp [0]),
    .X(\v0/z2/z1/q3 [1]));
 sky130_fd_sc_hd__and2_0 \v0/z2/z1/z4/z2/_0_  (.A(\v0/z2/z1/z4/temp [3]),
    .B(\v0/z2/z1/z4/temp [2]),
    .X(\v0/z2/z1/q3 [3]));
 sky130_fd_sc_hd__xor2_1 \v0/z2/z1/z4/z2/_1_  (.A(\v0/z2/z1/z4/temp [3]),
    .B(\v0/z2/z1/z4/temp [2]),
    .X(\v0/z2/z1/q3 [2]));
 sky130_fd_sc_hd__xnor2_1 \v0/z2/z1/z5/_07_  (.A(\v0/z2/z1/q0 [2]),
    .B(\v0/z2/z1/q1 [0]),
    .Y(\v0/z2/z1/z5/_00_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z2/z1/z5/_08_  (.A(\v0/z2/z1/_02_ ),
    .B(\v0/z2/z1/z5/_00_ ),
    .Y(\v0/z2/z1/q4 [0]));
 sky130_fd_sc_hd__maj3_1 \v0/z2/z1/z5/_09_  (.A(\v0/z2/z1/q0 [2]),
    .B(\v0/z2/z1/q1 [0]),
    .C(\v0/z2/z1/_02_ ),
    .X(\v0/z2/z1/z5/_01_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z2/z1/z5/_10_  (.A(\v0/z2/z1/q0 [3]),
    .B(\v0/z2/z1/q1 [1]),
    .Y(\v0/z2/z1/z5/_02_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z2/z1/z5/_11_  (.A(\v0/z2/z1/z5/_01_ ),
    .B(\v0/z2/z1/z5/_02_ ),
    .Y(\v0/z2/z1/q4 [1]));
 sky130_fd_sc_hd__maj3_1 \v0/z2/z1/z5/_12_  (.A(\v0/z2/z1/q0 [3]),
    .B(\v0/z2/z1/q1 [1]),
    .C(\v0/z2/z1/z5/_01_ ),
    .X(\v0/z2/z1/z5/_03_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z2/z1/z5/_13_  (.A(\v0/z2/z1/_00_ ),
    .B(\v0/z2/z1/q1 [2]),
    .Y(\v0/z2/z1/z5/_04_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z2/z1/z5/_14_  (.A(\v0/z2/z1/z5/_03_ ),
    .B(\v0/z2/z1/z5/_04_ ),
    .Y(\v0/z2/z1/q4 [2]));
 sky130_fd_sc_hd__maj3_1 \v0/z2/z1/z5/_15_  (.A(\v0/z2/z1/_00_ ),
    .B(\v0/z2/z1/q1 [2]),
    .C(\v0/z2/z1/z5/_03_ ),
    .X(\v0/z2/z1/z5/_05_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z2/z1/z5/_16_  (.A(\v0/z2/z1/_01_ ),
    .B(\v0/z2/z1/q1 [3]),
    .Y(\v0/z2/z1/z5/_06_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z2/z1/z5/_17_  (.A(\v0/z2/z1/z5/_05_ ),
    .B(\v0/z2/z1/z5/_06_ ),
    .Y(\v0/z2/z1/q4 [3]));
 sky130_fd_sc_hd__maj3_1 \v0/z2/z1/z5/_18_  (.A(\v0/z2/z1/_01_ ),
    .B(\v0/z2/z1/q1 [3]),
    .C(\v0/z2/z1/z5/_05_ ),
    .X(\v0/z2/z1/z5/Cout ));
 sky130_fd_sc_hd__xnor2_1 \v0/z2/z1/z6/_19_  (.A(\v0/z2/z1/_05_ ),
    .B(\v0/z2/z1/q2 [0]),
    .Y(\v0/z2/z1/z6/_00_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z2/z1/z6/_20_  (.A(\v0/z2/z1/_07_ ),
    .B(\v0/z2/z1/z6/_00_ ),
    .Y(\v0/z2/z1/q5 [0]));
 sky130_fd_sc_hd__maj3_1 \v0/z2/z1/z6/_21_  (.A(\v0/z2/z1/_05_ ),
    .B(\v0/z2/z1/q2 [0]),
    .C(\v0/z2/z1/_07_ ),
    .X(\v0/z2/z1/z6/_01_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z2/z1/z6/_22_  (.A(\v0/z2/z1/_06_ ),
    .B(\v0/z2/z1/q2 [1]),
    .Y(\v0/z2/z1/z6/_02_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z2/z1/z6/_23_  (.A(\v0/z2/z1/z6/_01_ ),
    .B(\v0/z2/z1/z6/_02_ ),
    .Y(\v0/z2/z1/q5 [1]));
 sky130_fd_sc_hd__maj3_1 \v0/z2/z1/z6/_24_  (.A(\v0/z2/z1/_06_ ),
    .B(\v0/z2/z1/q2 [1]),
    .C(\v0/z2/z1/z6/_01_ ),
    .X(\v0/z2/z1/z6/_03_ ));
 sky130_fd_sc_hd__lpflow_inputiso1p_1 \v0/z2/z1/z6/_25_  (.A(\v0/z2/z1/q3 [0]),
    .SLEEP(\v0/z2/z1/q2 [2]),
    .X(\v0/z2/z1/z6/_04_ ));
 sky130_fd_sc_hd__and2_0 \v0/z2/z1/z6/_26_  (.A(\v0/z2/z1/q3 [0]),
    .B(\v0/z2/z1/q2 [2]),
    .X(\v0/z2/z1/z6/_05_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z2/z1/z6/_27_  (.A(\v0/z2/z1/q3 [0]),
    .B(\v0/z2/z1/q2 [2]),
    .Y(\v0/z2/z1/z6/_06_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z2/z1/z6/_28_  (.A(\v0/z2/z1/z6/_04_ ),
    .B(\v0/z2/z1/z6/_06_ ),
    .Y(\v0/z2/z1/z6/_07_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z2/z1/z6/_29_  (.A(\v0/z2/z1/z6/_03_ ),
    .B(\v0/z2/z1/z6/_07_ ),
    .Y(\v0/z2/z1/q5 [2]));
 sky130_fd_sc_hd__nand2_1 \v0/z2/z1/z6/_30_  (.A(\v0/z2/z1/q3 [1]),
    .B(\v0/z2/z1/q2 [3]),
    .Y(\v0/z2/z1/z6/_08_ ));
 sky130_fd_sc_hd__xor2_1 \v0/z2/z1/z6/_31_  (.A(\v0/z2/z1/q3 [1]),
    .B(\v0/z2/z1/q2 [3]),
    .X(\v0/z2/z1/z6/_09_ ));
 sky130_fd_sc_hd__o21ai_0 \v0/z2/z1/z6/_32_  (.A1(\v0/z2/z1/z6/_03_ ),
    .A2(\v0/z2/z1/z6/_05_ ),
    .B1(\v0/z2/z1/z6/_04_ ),
    .Y(\v0/z2/z1/z6/_10_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z2/z1/z6/_33_  (.A(\v0/z2/z1/z6/_09_ ),
    .B(\v0/z2/z1/z6/_10_ ),
    .Y(\v0/z2/z1/q5 [3]));
 sky130_fd_sc_hd__nor2_1 \v0/z2/z1/z6/_34_  (.A(\v0/z2/z1/q3 [2]),
    .B(\v0/z2/z1/_03_ ),
    .Y(\v0/z2/z1/z6/_11_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z2/z1/z6/_35_  (.A(\v0/z2/z1/q3 [2]),
    .B(\v0/z2/z1/_03_ ),
    .Y(\v0/z2/z1/z6/_12_ ));
 sky130_fd_sc_hd__nand2b_1 \v0/z2/z1/z6/_36_  (.A_N(\v0/z2/z1/z6/_11_ ),
    .B(\v0/z2/z1/z6/_12_ ),
    .Y(\v0/z2/z1/z6/_13_ ));
 sky130_fd_sc_hd__o221ai_1 \v0/z2/z1/z6/_37_  (.A1(\v0/z2/z1/q3 [1]),
    .A2(\v0/z2/z1/q2 [3]),
    .B1(\v0/z2/z1/z6/_03_ ),
    .B2(\v0/z2/z1/z6/_05_ ),
    .C1(\v0/z2/z1/z6/_04_ ),
    .Y(\v0/z2/z1/z6/_14_ ));
 sky130_fd_sc_hd__a21oi_1 \v0/z2/z1/z6/_38_  (.A1(\v0/z2/z1/z6/_08_ ),
    .A2(\v0/z2/z1/z6/_14_ ),
    .B1(\v0/z2/z1/z6/_13_ ),
    .Y(\v0/z2/z1/z6/_15_ ));
 sky130_fd_sc_hd__and3_1 \v0/z2/z1/z6/_39_  (.A(\v0/z2/z1/z6/_08_ ),
    .B(\v0/z2/z1/z6/_13_ ),
    .C(\v0/z2/z1/z6/_14_ ),
    .X(\v0/z2/z1/z6/_16_ ));
 sky130_fd_sc_hd__nor2_1 \v0/z2/z1/z6/_40_  (.A(\v0/z2/z1/z6/_15_ ),
    .B(\v0/z2/z1/z6/_16_ ),
    .Y(\v0/z2/z1/q5 [4]));
 sky130_fd_sc_hd__xnor2_1 \v0/z2/z1/z6/_41_  (.A(\v0/z2/z1/q3 [3]),
    .B(\v0/z2/z1/_04_ ),
    .Y(\v0/z2/z1/z6/_17_ ));
 sky130_fd_sc_hd__a31oi_1 \v0/z2/z1/z6/_42_  (.A1(\v0/z2/z1/z6/_08_ ),
    .A2(\v0/z2/z1/z6/_12_ ),
    .A3(\v0/z2/z1/z6/_14_ ),
    .B1(\v0/z2/z1/z6/_11_ ),
    .Y(\v0/z2/z1/z6/_18_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z2/z1/z6/_43_  (.A(\v0/z2/z1/z6/_17_ ),
    .B(\v0/z2/z1/z6/_18_ ),
    .Y(\v0/z2/z1/q5 [5]));
 sky130_fd_sc_hd__maj3_1 \v0/z2/z1/z6/_44_  (.A(\v0/z2/z1/q3 [3]),
    .B(\v0/z2/z1/_04_ ),
    .C(\v0/z2/z1/z6/_18_ ),
    .X(\v0/z2/z1/z6/Cout ));
 sky130_fd_sc_hd__xnor2_1 \v0/z2/z1/z7/_19_  (.A(\v0/z2/z1/q5 [0]),
    .B(\v0/z2/z1/q4 [0]),
    .Y(\v0/z2/z1/z7/_00_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z2/z1/z7/_20_  (.A(\v0/z2/z1/_10_ ),
    .B(\v0/z2/z1/z7/_00_ ),
    .Y(\v0/q1 [2]));
 sky130_fd_sc_hd__maj3_1 \v0/z2/z1/z7/_21_  (.A(\v0/z2/z1/q5 [0]),
    .B(\v0/z2/z1/q4 [0]),
    .C(\v0/z2/z1/_10_ ),
    .X(\v0/z2/z1/z7/_01_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z2/z1/z7/_22_  (.A(\v0/z2/z1/q5 [1]),
    .B(\v0/z2/z1/q4 [1]),
    .Y(\v0/z2/z1/z7/_02_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z2/z1/z7/_23_  (.A(\v0/z2/z1/z7/_01_ ),
    .B(\v0/z2/z1/z7/_02_ ),
    .Y(\v0/q1 [3]));
 sky130_fd_sc_hd__maj3_1 \v0/z2/z1/z7/_24_  (.A(\v0/z2/z1/q5 [1]),
    .B(\v0/z2/z1/q4 [1]),
    .C(\v0/z2/z1/z7/_01_ ),
    .X(\v0/z2/z1/z7/_03_ ));
 sky130_fd_sc_hd__lpflow_inputiso1p_1 \v0/z2/z1/z7/_25_  (.A(\v0/z2/z1/q5 [2]),
    .SLEEP(\v0/z2/z1/q4 [2]),
    .X(\v0/z2/z1/z7/_04_ ));
 sky130_fd_sc_hd__and2_0 \v0/z2/z1/z7/_26_  (.A(\v0/z2/z1/q5 [2]),
    .B(\v0/z2/z1/q4 [2]),
    .X(\v0/z2/z1/z7/_05_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z2/z1/z7/_27_  (.A(\v0/z2/z1/q5 [2]),
    .B(\v0/z2/z1/q4 [2]),
    .Y(\v0/z2/z1/z7/_06_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z2/z1/z7/_28_  (.A(\v0/z2/z1/z7/_04_ ),
    .B(\v0/z2/z1/z7/_06_ ),
    .Y(\v0/z2/z1/z7/_07_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z2/z1/z7/_29_  (.A(\v0/z2/z1/z7/_03_ ),
    .B(\v0/z2/z1/z7/_07_ ),
    .Y(\v0/z2/q0 [4]));
 sky130_fd_sc_hd__nand2_1 \v0/z2/z1/z7/_30_  (.A(\v0/z2/z1/q5 [3]),
    .B(\v0/z2/z1/q4 [3]),
    .Y(\v0/z2/z1/z7/_08_ ));
 sky130_fd_sc_hd__xor2_1 \v0/z2/z1/z7/_31_  (.A(\v0/z2/z1/q5 [3]),
    .B(\v0/z2/z1/q4 [3]),
    .X(\v0/z2/z1/z7/_09_ ));
 sky130_fd_sc_hd__o21ai_0 \v0/z2/z1/z7/_32_  (.A1(\v0/z2/z1/z7/_03_ ),
    .A2(\v0/z2/z1/z7/_05_ ),
    .B1(\v0/z2/z1/z7/_04_ ),
    .Y(\v0/z2/z1/z7/_10_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z2/z1/z7/_33_  (.A(\v0/z2/z1/z7/_09_ ),
    .B(\v0/z2/z1/z7/_10_ ),
    .Y(\v0/z2/q0 [5]));
 sky130_fd_sc_hd__nor2_1 \v0/z2/z1/z7/_34_  (.A(\v0/z2/z1/q5 [4]),
    .B(\v0/z2/z1/_08_ ),
    .Y(\v0/z2/z1/z7/_11_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z2/z1/z7/_35_  (.A(\v0/z2/z1/q5 [4]),
    .B(\v0/z2/z1/_08_ ),
    .Y(\v0/z2/z1/z7/_12_ ));
 sky130_fd_sc_hd__nand2b_1 \v0/z2/z1/z7/_36_  (.A_N(\v0/z2/z1/z7/_11_ ),
    .B(\v0/z2/z1/z7/_12_ ),
    .Y(\v0/z2/z1/z7/_13_ ));
 sky130_fd_sc_hd__o221ai_1 \v0/z2/z1/z7/_37_  (.A1(\v0/z2/z1/q5 [3]),
    .A2(\v0/z2/z1/q4 [3]),
    .B1(\v0/z2/z1/z7/_03_ ),
    .B2(\v0/z2/z1/z7/_05_ ),
    .C1(\v0/z2/z1/z7/_04_ ),
    .Y(\v0/z2/z1/z7/_14_ ));
 sky130_fd_sc_hd__a21oi_1 \v0/z2/z1/z7/_38_  (.A1(\v0/z2/z1/z7/_08_ ),
    .A2(\v0/z2/z1/z7/_14_ ),
    .B1(\v0/z2/z1/z7/_13_ ),
    .Y(\v0/z2/z1/z7/_15_ ));
 sky130_fd_sc_hd__and3_1 \v0/z2/z1/z7/_39_  (.A(\v0/z2/z1/z7/_08_ ),
    .B(\v0/z2/z1/z7/_13_ ),
    .C(\v0/z2/z1/z7/_14_ ),
    .X(\v0/z2/z1/z7/_16_ ));
 sky130_fd_sc_hd__nor2_1 \v0/z2/z1/z7/_40_  (.A(\v0/z2/z1/z7/_15_ ),
    .B(\v0/z2/z1/z7/_16_ ),
    .Y(\v0/z2/q0 [6]));
 sky130_fd_sc_hd__xnor2_1 \v0/z2/z1/z7/_41_  (.A(\v0/z2/z1/q5 [5]),
    .B(\v0/z2/z1/_09_ ),
    .Y(\v0/z2/z1/z7/_17_ ));
 sky130_fd_sc_hd__a31oi_1 \v0/z2/z1/z7/_42_  (.A1(\v0/z2/z1/z7/_08_ ),
    .A2(\v0/z2/z1/z7/_12_ ),
    .A3(\v0/z2/z1/z7/_14_ ),
    .B1(\v0/z2/z1/z7/_11_ ),
    .Y(\v0/z2/z1/z7/_18_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z2/z1/z7/_43_  (.A(\v0/z2/z1/z7/_17_ ),
    .B(\v0/z2/z1/z7/_18_ ),
    .Y(\v0/z2/q0 [7]));
 sky130_fd_sc_hd__maj3_1 \v0/z2/z1/z7/_44_  (.A(\v0/z2/z1/q5 [5]),
    .B(\v0/z2/z1/_09_ ),
    .C(\v0/z2/z1/z7/_18_ ),
    .X(\v0/z2/z1/z7/Cout ));
 sky130_fd_sc_hd__conb_1 \v0/z2/z2/_11_  (.LO(\v0/z2/z2/_00_ ));
 sky130_fd_sc_hd__conb_1 \v0/z2/z2/_12_  (.LO(\v0/z2/z2/_01_ ));
 sky130_fd_sc_hd__conb_1 \v0/z2/z2/_13_  (.LO(\v0/z2/z2/_02_ ));
 sky130_fd_sc_hd__conb_1 \v0/z2/z2/_14_  (.LO(\v0/z2/z2/_03_ ));
 sky130_fd_sc_hd__conb_1 \v0/z2/z2/_15_  (.LO(\v0/z2/z2/_04_ ));
 sky130_fd_sc_hd__conb_1 \v0/z2/z2/_16_  (.LO(\v0/z2/z2/_05_ ));
 sky130_fd_sc_hd__conb_1 \v0/z2/z2/_17_  (.LO(\v0/z2/z2/_06_ ));
 sky130_fd_sc_hd__conb_1 \v0/z2/z2/_18_  (.LO(\v0/z2/z2/_07_ ));
 sky130_fd_sc_hd__conb_1 \v0/z2/z2/_19_  (.LO(\v0/z2/z2/_08_ ));
 sky130_fd_sc_hd__conb_1 \v0/z2/z2/_20_  (.LO(\v0/z2/z2/_09_ ));
 sky130_fd_sc_hd__conb_1 \v0/z2/z2/_21_  (.LO(\v0/z2/z2/_10_ ));
 sky130_fd_sc_hd__and2_0 \v0/z2/z2/z1/_0_  (.A(b[0]),
    .B(abs_a[12]),
    .X(\v0/z2/q1 [0]));
 sky130_fd_sc_hd__and2_0 \v0/z2/z2/z1/_1_  (.A(b[0]),
    .B(abs_a[13]),
    .X(\v0/z2/z2/z1/temp [0]));
 sky130_fd_sc_hd__and2_0 \v0/z2/z2/z1/_2_  (.A(abs_a[12]),
    .B(abs_b[1]),
    .X(\v0/z2/z2/z1/temp [1]));
 sky130_fd_sc_hd__and2_0 \v0/z2/z2/z1/_3_  (.A(abs_a[13]),
    .B(abs_b[1]),
    .X(\v0/z2/z2/z1/temp [2]));
 sky130_fd_sc_hd__and2_0 \v0/z2/z2/z1/z1/_0_  (.A(\v0/z2/z2/z1/temp [1]),
    .B(\v0/z2/z2/z1/temp [0]),
    .X(\v0/z2/z2/z1/temp [3]));
 sky130_fd_sc_hd__xor2_1 \v0/z2/z2/z1/z1/_1_  (.A(\v0/z2/z2/z1/temp [1]),
    .B(\v0/z2/z2/z1/temp [0]),
    .X(\v0/z2/q1 [1]));
 sky130_fd_sc_hd__and2_0 \v0/z2/z2/z1/z2/_0_  (.A(\v0/z2/z2/z1/temp [3]),
    .B(\v0/z2/z2/z1/temp [2]),
    .X(\v0/z2/z2/q0 [3]));
 sky130_fd_sc_hd__xor2_1 \v0/z2/z2/z1/z2/_1_  (.A(\v0/z2/z2/z1/temp [3]),
    .B(\v0/z2/z2/z1/temp [2]),
    .X(\v0/z2/z2/q0 [2]));
 sky130_fd_sc_hd__and2_0 \v0/z2/z2/z2/_0_  (.A(b[0]),
    .B(abs_a[14]),
    .X(\v0/z2/z2/q1 [0]));
 sky130_fd_sc_hd__and2_0 \v0/z2/z2/z2/_1_  (.A(b[0]),
    .B(abs_a[15]),
    .X(\v0/z2/z2/z2/temp [0]));
 sky130_fd_sc_hd__and2_0 \v0/z2/z2/z2/_2_  (.A(abs_a[14]),
    .B(abs_b[1]),
    .X(\v0/z2/z2/z2/temp [1]));
 sky130_fd_sc_hd__and2_0 \v0/z2/z2/z2/_3_  (.A(abs_a[15]),
    .B(abs_b[1]),
    .X(\v0/z2/z2/z2/temp [2]));
 sky130_fd_sc_hd__and2_0 \v0/z2/z2/z2/z1/_0_  (.A(\v0/z2/z2/z2/temp [1]),
    .B(\v0/z2/z2/z2/temp [0]),
    .X(\v0/z2/z2/z2/temp [3]));
 sky130_fd_sc_hd__xor2_1 \v0/z2/z2/z2/z1/_1_  (.A(\v0/z2/z2/z2/temp [1]),
    .B(\v0/z2/z2/z2/temp [0]),
    .X(\v0/z2/z2/q1 [1]));
 sky130_fd_sc_hd__and2_0 \v0/z2/z2/z2/z2/_0_  (.A(\v0/z2/z2/z2/temp [3]),
    .B(\v0/z2/z2/z2/temp [2]),
    .X(\v0/z2/z2/q1 [3]));
 sky130_fd_sc_hd__xor2_1 \v0/z2/z2/z2/z2/_1_  (.A(\v0/z2/z2/z2/temp [3]),
    .B(\v0/z2/z2/z2/temp [2]),
    .X(\v0/z2/z2/q1 [2]));
 sky130_fd_sc_hd__and2_0 \v0/z2/z2/z3/_0_  (.A(abs_b[2]),
    .B(abs_a[12]),
    .X(\v0/z2/z2/q2 [0]));
 sky130_fd_sc_hd__and2_0 \v0/z2/z2/z3/_1_  (.A(abs_b[2]),
    .B(abs_a[13]),
    .X(\v0/z2/z2/z3/temp [0]));
 sky130_fd_sc_hd__and2_0 \v0/z2/z2/z3/_2_  (.A(abs_a[12]),
    .B(abs_b[3]),
    .X(\v0/z2/z2/z3/temp [1]));
 sky130_fd_sc_hd__and2_0 \v0/z2/z2/z3/_3_  (.A(abs_a[13]),
    .B(abs_b[3]),
    .X(\v0/z2/z2/z3/temp [2]));
 sky130_fd_sc_hd__and2_0 \v0/z2/z2/z3/z1/_0_  (.A(\v0/z2/z2/z3/temp [1]),
    .B(\v0/z2/z2/z3/temp [0]),
    .X(\v0/z2/z2/z3/temp [3]));
 sky130_fd_sc_hd__xor2_1 \v0/z2/z2/z3/z1/_1_  (.A(\v0/z2/z2/z3/temp [1]),
    .B(\v0/z2/z2/z3/temp [0]),
    .X(\v0/z2/z2/q2 [1]));
 sky130_fd_sc_hd__and2_0 \v0/z2/z2/z3/z2/_0_  (.A(\v0/z2/z2/z3/temp [3]),
    .B(\v0/z2/z2/z3/temp [2]),
    .X(\v0/z2/z2/q2 [3]));
 sky130_fd_sc_hd__xor2_1 \v0/z2/z2/z3/z2/_1_  (.A(\v0/z2/z2/z3/temp [3]),
    .B(\v0/z2/z2/z3/temp [2]),
    .X(\v0/z2/z2/q2 [2]));
 sky130_fd_sc_hd__and2_0 \v0/z2/z2/z4/_0_  (.A(abs_b[2]),
    .B(abs_a[14]),
    .X(\v0/z2/z2/q3 [0]));
 sky130_fd_sc_hd__and2_0 \v0/z2/z2/z4/_1_  (.A(abs_b[2]),
    .B(abs_a[15]),
    .X(\v0/z2/z2/z4/temp [0]));
 sky130_fd_sc_hd__and2_0 \v0/z2/z2/z4/_2_  (.A(abs_a[14]),
    .B(abs_b[3]),
    .X(\v0/z2/z2/z4/temp [1]));
 sky130_fd_sc_hd__and2_0 \v0/z2/z2/z4/_3_  (.A(abs_a[15]),
    .B(abs_b[3]),
    .X(\v0/z2/z2/z4/temp [2]));
 sky130_fd_sc_hd__and2_0 \v0/z2/z2/z4/z1/_0_  (.A(\v0/z2/z2/z4/temp [1]),
    .B(\v0/z2/z2/z4/temp [0]),
    .X(\v0/z2/z2/z4/temp [3]));
 sky130_fd_sc_hd__xor2_1 \v0/z2/z2/z4/z1/_1_  (.A(\v0/z2/z2/z4/temp [1]),
    .B(\v0/z2/z2/z4/temp [0]),
    .X(\v0/z2/z2/q3 [1]));
 sky130_fd_sc_hd__and2_0 \v0/z2/z2/z4/z2/_0_  (.A(\v0/z2/z2/z4/temp [3]),
    .B(\v0/z2/z2/z4/temp [2]),
    .X(\v0/z2/z2/q3 [3]));
 sky130_fd_sc_hd__xor2_1 \v0/z2/z2/z4/z2/_1_  (.A(\v0/z2/z2/z4/temp [3]),
    .B(\v0/z2/z2/z4/temp [2]),
    .X(\v0/z2/z2/q3 [2]));
 sky130_fd_sc_hd__xnor2_1 \v0/z2/z2/z5/_07_  (.A(\v0/z2/z2/q0 [2]),
    .B(\v0/z2/z2/q1 [0]),
    .Y(\v0/z2/z2/z5/_00_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z2/z2/z5/_08_  (.A(\v0/z2/z2/_02_ ),
    .B(\v0/z2/z2/z5/_00_ ),
    .Y(\v0/z2/z2/q4 [0]));
 sky130_fd_sc_hd__maj3_1 \v0/z2/z2/z5/_09_  (.A(\v0/z2/z2/q0 [2]),
    .B(\v0/z2/z2/q1 [0]),
    .C(\v0/z2/z2/_02_ ),
    .X(\v0/z2/z2/z5/_01_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z2/z2/z5/_10_  (.A(\v0/z2/z2/q0 [3]),
    .B(\v0/z2/z2/q1 [1]),
    .Y(\v0/z2/z2/z5/_02_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z2/z2/z5/_11_  (.A(\v0/z2/z2/z5/_01_ ),
    .B(\v0/z2/z2/z5/_02_ ),
    .Y(\v0/z2/z2/q4 [1]));
 sky130_fd_sc_hd__maj3_1 \v0/z2/z2/z5/_12_  (.A(\v0/z2/z2/q0 [3]),
    .B(\v0/z2/z2/q1 [1]),
    .C(\v0/z2/z2/z5/_01_ ),
    .X(\v0/z2/z2/z5/_03_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z2/z2/z5/_13_  (.A(\v0/z2/z2/_00_ ),
    .B(\v0/z2/z2/q1 [2]),
    .Y(\v0/z2/z2/z5/_04_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z2/z2/z5/_14_  (.A(\v0/z2/z2/z5/_03_ ),
    .B(\v0/z2/z2/z5/_04_ ),
    .Y(\v0/z2/z2/q4 [2]));
 sky130_fd_sc_hd__maj3_1 \v0/z2/z2/z5/_15_  (.A(\v0/z2/z2/_00_ ),
    .B(\v0/z2/z2/q1 [2]),
    .C(\v0/z2/z2/z5/_03_ ),
    .X(\v0/z2/z2/z5/_05_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z2/z2/z5/_16_  (.A(\v0/z2/z2/_01_ ),
    .B(\v0/z2/z2/q1 [3]),
    .Y(\v0/z2/z2/z5/_06_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z2/z2/z5/_17_  (.A(\v0/z2/z2/z5/_05_ ),
    .B(\v0/z2/z2/z5/_06_ ),
    .Y(\v0/z2/z2/q4 [3]));
 sky130_fd_sc_hd__maj3_1 \v0/z2/z2/z5/_18_  (.A(\v0/z2/z2/_01_ ),
    .B(\v0/z2/z2/q1 [3]),
    .C(\v0/z2/z2/z5/_05_ ),
    .X(\v0/z2/z2/z5/Cout ));
 sky130_fd_sc_hd__xnor2_1 \v0/z2/z2/z6/_19_  (.A(\v0/z2/z2/_05_ ),
    .B(\v0/z2/z2/q2 [0]),
    .Y(\v0/z2/z2/z6/_00_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z2/z2/z6/_20_  (.A(\v0/z2/z2/_07_ ),
    .B(\v0/z2/z2/z6/_00_ ),
    .Y(\v0/z2/z2/q5 [0]));
 sky130_fd_sc_hd__maj3_1 \v0/z2/z2/z6/_21_  (.A(\v0/z2/z2/_05_ ),
    .B(\v0/z2/z2/q2 [0]),
    .C(\v0/z2/z2/_07_ ),
    .X(\v0/z2/z2/z6/_01_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z2/z2/z6/_22_  (.A(\v0/z2/z2/_06_ ),
    .B(\v0/z2/z2/q2 [1]),
    .Y(\v0/z2/z2/z6/_02_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z2/z2/z6/_23_  (.A(\v0/z2/z2/z6/_01_ ),
    .B(\v0/z2/z2/z6/_02_ ),
    .Y(\v0/z2/z2/q5 [1]));
 sky130_fd_sc_hd__maj3_1 \v0/z2/z2/z6/_24_  (.A(\v0/z2/z2/_06_ ),
    .B(\v0/z2/z2/q2 [1]),
    .C(\v0/z2/z2/z6/_01_ ),
    .X(\v0/z2/z2/z6/_03_ ));
 sky130_fd_sc_hd__lpflow_inputiso1p_1 \v0/z2/z2/z6/_25_  (.A(\v0/z2/z2/q3 [0]),
    .SLEEP(\v0/z2/z2/q2 [2]),
    .X(\v0/z2/z2/z6/_04_ ));
 sky130_fd_sc_hd__and2_0 \v0/z2/z2/z6/_26_  (.A(\v0/z2/z2/q3 [0]),
    .B(\v0/z2/z2/q2 [2]),
    .X(\v0/z2/z2/z6/_05_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z2/z2/z6/_27_  (.A(\v0/z2/z2/q3 [0]),
    .B(\v0/z2/z2/q2 [2]),
    .Y(\v0/z2/z2/z6/_06_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z2/z2/z6/_28_  (.A(\v0/z2/z2/z6/_04_ ),
    .B(\v0/z2/z2/z6/_06_ ),
    .Y(\v0/z2/z2/z6/_07_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z2/z2/z6/_29_  (.A(\v0/z2/z2/z6/_03_ ),
    .B(\v0/z2/z2/z6/_07_ ),
    .Y(\v0/z2/z2/q5 [2]));
 sky130_fd_sc_hd__nand2_1 \v0/z2/z2/z6/_30_  (.A(\v0/z2/z2/q3 [1]),
    .B(\v0/z2/z2/q2 [3]),
    .Y(\v0/z2/z2/z6/_08_ ));
 sky130_fd_sc_hd__xor2_1 \v0/z2/z2/z6/_31_  (.A(\v0/z2/z2/q3 [1]),
    .B(\v0/z2/z2/q2 [3]),
    .X(\v0/z2/z2/z6/_09_ ));
 sky130_fd_sc_hd__o21ai_0 \v0/z2/z2/z6/_32_  (.A1(\v0/z2/z2/z6/_03_ ),
    .A2(\v0/z2/z2/z6/_05_ ),
    .B1(\v0/z2/z2/z6/_04_ ),
    .Y(\v0/z2/z2/z6/_10_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z2/z2/z6/_33_  (.A(\v0/z2/z2/z6/_09_ ),
    .B(\v0/z2/z2/z6/_10_ ),
    .Y(\v0/z2/z2/q5 [3]));
 sky130_fd_sc_hd__nor2_1 \v0/z2/z2/z6/_34_  (.A(\v0/z2/z2/q3 [2]),
    .B(\v0/z2/z2/_03_ ),
    .Y(\v0/z2/z2/z6/_11_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z2/z2/z6/_35_  (.A(\v0/z2/z2/q3 [2]),
    .B(\v0/z2/z2/_03_ ),
    .Y(\v0/z2/z2/z6/_12_ ));
 sky130_fd_sc_hd__nand2b_1 \v0/z2/z2/z6/_36_  (.A_N(\v0/z2/z2/z6/_11_ ),
    .B(\v0/z2/z2/z6/_12_ ),
    .Y(\v0/z2/z2/z6/_13_ ));
 sky130_fd_sc_hd__o221ai_1 \v0/z2/z2/z6/_37_  (.A1(\v0/z2/z2/q3 [1]),
    .A2(\v0/z2/z2/q2 [3]),
    .B1(\v0/z2/z2/z6/_03_ ),
    .B2(\v0/z2/z2/z6/_05_ ),
    .C1(\v0/z2/z2/z6/_04_ ),
    .Y(\v0/z2/z2/z6/_14_ ));
 sky130_fd_sc_hd__a21oi_1 \v0/z2/z2/z6/_38_  (.A1(\v0/z2/z2/z6/_08_ ),
    .A2(\v0/z2/z2/z6/_14_ ),
    .B1(\v0/z2/z2/z6/_13_ ),
    .Y(\v0/z2/z2/z6/_15_ ));
 sky130_fd_sc_hd__and3_1 \v0/z2/z2/z6/_39_  (.A(\v0/z2/z2/z6/_08_ ),
    .B(\v0/z2/z2/z6/_13_ ),
    .C(\v0/z2/z2/z6/_14_ ),
    .X(\v0/z2/z2/z6/_16_ ));
 sky130_fd_sc_hd__nor2_1 \v0/z2/z2/z6/_40_  (.A(\v0/z2/z2/z6/_15_ ),
    .B(\v0/z2/z2/z6/_16_ ),
    .Y(\v0/z2/z2/q5 [4]));
 sky130_fd_sc_hd__xnor2_1 \v0/z2/z2/z6/_41_  (.A(\v0/z2/z2/q3 [3]),
    .B(\v0/z2/z2/_04_ ),
    .Y(\v0/z2/z2/z6/_17_ ));
 sky130_fd_sc_hd__a31oi_1 \v0/z2/z2/z6/_42_  (.A1(\v0/z2/z2/z6/_08_ ),
    .A2(\v0/z2/z2/z6/_12_ ),
    .A3(\v0/z2/z2/z6/_14_ ),
    .B1(\v0/z2/z2/z6/_11_ ),
    .Y(\v0/z2/z2/z6/_18_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z2/z2/z6/_43_  (.A(\v0/z2/z2/z6/_17_ ),
    .B(\v0/z2/z2/z6/_18_ ),
    .Y(\v0/z2/z2/q5 [5]));
 sky130_fd_sc_hd__maj3_1 \v0/z2/z2/z6/_44_  (.A(\v0/z2/z2/q3 [3]),
    .B(\v0/z2/z2/_04_ ),
    .C(\v0/z2/z2/z6/_18_ ),
    .X(\v0/z2/z2/z6/Cout ));
 sky130_fd_sc_hd__xnor2_1 \v0/z2/z2/z7/_19_  (.A(\v0/z2/z2/q5 [0]),
    .B(\v0/z2/z2/q4 [0]),
    .Y(\v0/z2/z2/z7/_00_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z2/z2/z7/_20_  (.A(\v0/z2/z2/_10_ ),
    .B(\v0/z2/z2/z7/_00_ ),
    .Y(\v0/z2/q1 [2]));
 sky130_fd_sc_hd__maj3_1 \v0/z2/z2/z7/_21_  (.A(\v0/z2/z2/q5 [0]),
    .B(\v0/z2/z2/q4 [0]),
    .C(\v0/z2/z2/_10_ ),
    .X(\v0/z2/z2/z7/_01_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z2/z2/z7/_22_  (.A(\v0/z2/z2/q5 [1]),
    .B(\v0/z2/z2/q4 [1]),
    .Y(\v0/z2/z2/z7/_02_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z2/z2/z7/_23_  (.A(\v0/z2/z2/z7/_01_ ),
    .B(\v0/z2/z2/z7/_02_ ),
    .Y(\v0/z2/q1 [3]));
 sky130_fd_sc_hd__maj3_1 \v0/z2/z2/z7/_24_  (.A(\v0/z2/z2/q5 [1]),
    .B(\v0/z2/z2/q4 [1]),
    .C(\v0/z2/z2/z7/_01_ ),
    .X(\v0/z2/z2/z7/_03_ ));
 sky130_fd_sc_hd__lpflow_inputiso1p_1 \v0/z2/z2/z7/_25_  (.A(\v0/z2/z2/q5 [2]),
    .SLEEP(\v0/z2/z2/q4 [2]),
    .X(\v0/z2/z2/z7/_04_ ));
 sky130_fd_sc_hd__and2_0 \v0/z2/z2/z7/_26_  (.A(\v0/z2/z2/q5 [2]),
    .B(\v0/z2/z2/q4 [2]),
    .X(\v0/z2/z2/z7/_05_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z2/z2/z7/_27_  (.A(\v0/z2/z2/q5 [2]),
    .B(\v0/z2/z2/q4 [2]),
    .Y(\v0/z2/z2/z7/_06_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z2/z2/z7/_28_  (.A(\v0/z2/z2/z7/_04_ ),
    .B(\v0/z2/z2/z7/_06_ ),
    .Y(\v0/z2/z2/z7/_07_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z2/z2/z7/_29_  (.A(\v0/z2/z2/z7/_03_ ),
    .B(\v0/z2/z2/z7/_07_ ),
    .Y(\v0/z2/q1 [4]));
 sky130_fd_sc_hd__nand2_1 \v0/z2/z2/z7/_30_  (.A(\v0/z2/z2/q5 [3]),
    .B(\v0/z2/z2/q4 [3]),
    .Y(\v0/z2/z2/z7/_08_ ));
 sky130_fd_sc_hd__xor2_1 \v0/z2/z2/z7/_31_  (.A(\v0/z2/z2/q5 [3]),
    .B(\v0/z2/z2/q4 [3]),
    .X(\v0/z2/z2/z7/_09_ ));
 sky130_fd_sc_hd__o21ai_0 \v0/z2/z2/z7/_32_  (.A1(\v0/z2/z2/z7/_03_ ),
    .A2(\v0/z2/z2/z7/_05_ ),
    .B1(\v0/z2/z2/z7/_04_ ),
    .Y(\v0/z2/z2/z7/_10_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z2/z2/z7/_33_  (.A(\v0/z2/z2/z7/_09_ ),
    .B(\v0/z2/z2/z7/_10_ ),
    .Y(\v0/z2/q1 [5]));
 sky130_fd_sc_hd__nor2_1 \v0/z2/z2/z7/_34_  (.A(\v0/z2/z2/q5 [4]),
    .B(\v0/z2/z2/_08_ ),
    .Y(\v0/z2/z2/z7/_11_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z2/z2/z7/_35_  (.A(\v0/z2/z2/q5 [4]),
    .B(\v0/z2/z2/_08_ ),
    .Y(\v0/z2/z2/z7/_12_ ));
 sky130_fd_sc_hd__nand2b_1 \v0/z2/z2/z7/_36_  (.A_N(\v0/z2/z2/z7/_11_ ),
    .B(\v0/z2/z2/z7/_12_ ),
    .Y(\v0/z2/z2/z7/_13_ ));
 sky130_fd_sc_hd__o221ai_1 \v0/z2/z2/z7/_37_  (.A1(\v0/z2/z2/q5 [3]),
    .A2(\v0/z2/z2/q4 [3]),
    .B1(\v0/z2/z2/z7/_03_ ),
    .B2(\v0/z2/z2/z7/_05_ ),
    .C1(\v0/z2/z2/z7/_04_ ),
    .Y(\v0/z2/z2/z7/_14_ ));
 sky130_fd_sc_hd__a21oi_1 \v0/z2/z2/z7/_38_  (.A1(\v0/z2/z2/z7/_08_ ),
    .A2(\v0/z2/z2/z7/_14_ ),
    .B1(\v0/z2/z2/z7/_13_ ),
    .Y(\v0/z2/z2/z7/_15_ ));
 sky130_fd_sc_hd__and3_1 \v0/z2/z2/z7/_39_  (.A(\v0/z2/z2/z7/_08_ ),
    .B(\v0/z2/z2/z7/_13_ ),
    .C(\v0/z2/z2/z7/_14_ ),
    .X(\v0/z2/z2/z7/_16_ ));
 sky130_fd_sc_hd__nor2_1 \v0/z2/z2/z7/_40_  (.A(\v0/z2/z2/z7/_15_ ),
    .B(\v0/z2/z2/z7/_16_ ),
    .Y(\v0/z2/q1 [6]));
 sky130_fd_sc_hd__xnor2_1 \v0/z2/z2/z7/_41_  (.A(\v0/z2/z2/q5 [5]),
    .B(\v0/z2/z2/_09_ ),
    .Y(\v0/z2/z2/z7/_17_ ));
 sky130_fd_sc_hd__a31oi_1 \v0/z2/z2/z7/_42_  (.A1(\v0/z2/z2/z7/_08_ ),
    .A2(\v0/z2/z2/z7/_12_ ),
    .A3(\v0/z2/z2/z7/_14_ ),
    .B1(\v0/z2/z2/z7/_11_ ),
    .Y(\v0/z2/z2/z7/_18_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z2/z2/z7/_43_  (.A(\v0/z2/z2/z7/_17_ ),
    .B(\v0/z2/z2/z7/_18_ ),
    .Y(\v0/z2/q1 [7]));
 sky130_fd_sc_hd__maj3_1 \v0/z2/z2/z7/_44_  (.A(\v0/z2/z2/q5 [5]),
    .B(\v0/z2/z2/_09_ ),
    .C(\v0/z2/z2/z7/_18_ ),
    .X(\v0/z2/z2/z7/Cout ));
 sky130_fd_sc_hd__conb_1 \v0/z2/z3/_11_  (.LO(\v0/z2/z3/_00_ ));
 sky130_fd_sc_hd__conb_1 \v0/z2/z3/_12_  (.LO(\v0/z2/z3/_01_ ));
 sky130_fd_sc_hd__conb_1 \v0/z2/z3/_13_  (.LO(\v0/z2/z3/_02_ ));
 sky130_fd_sc_hd__conb_1 \v0/z2/z3/_14_  (.LO(\v0/z2/z3/_03_ ));
 sky130_fd_sc_hd__conb_1 \v0/z2/z3/_15_  (.LO(\v0/z2/z3/_04_ ));
 sky130_fd_sc_hd__conb_1 \v0/z2/z3/_16_  (.LO(\v0/z2/z3/_05_ ));
 sky130_fd_sc_hd__conb_1 \v0/z2/z3/_17_  (.LO(\v0/z2/z3/_06_ ));
 sky130_fd_sc_hd__conb_1 \v0/z2/z3/_18_  (.LO(\v0/z2/z3/_07_ ));
 sky130_fd_sc_hd__conb_1 \v0/z2/z3/_19_  (.LO(\v0/z2/z3/_08_ ));
 sky130_fd_sc_hd__conb_1 \v0/z2/z3/_20_  (.LO(\v0/z2/z3/_09_ ));
 sky130_fd_sc_hd__conb_1 \v0/z2/z3/_21_  (.LO(\v0/z2/z3/_10_ ));
 sky130_fd_sc_hd__and2_0 \v0/z2/z3/z1/_0_  (.A(abs_b[4]),
    .B(abs_a[8]),
    .X(\v0/z2/q2 [0]));
 sky130_fd_sc_hd__and2_0 \v0/z2/z3/z1/_1_  (.A(abs_b[4]),
    .B(abs_a[9]),
    .X(\v0/z2/z3/z1/temp [0]));
 sky130_fd_sc_hd__and2_0 \v0/z2/z3/z1/_2_  (.A(abs_a[8]),
    .B(abs_b[5]),
    .X(\v0/z2/z3/z1/temp [1]));
 sky130_fd_sc_hd__and2_0 \v0/z2/z3/z1/_3_  (.A(abs_a[9]),
    .B(abs_b[5]),
    .X(\v0/z2/z3/z1/temp [2]));
 sky130_fd_sc_hd__and2_0 \v0/z2/z3/z1/z1/_0_  (.A(\v0/z2/z3/z1/temp [1]),
    .B(\v0/z2/z3/z1/temp [0]),
    .X(\v0/z2/z3/z1/temp [3]));
 sky130_fd_sc_hd__xor2_1 \v0/z2/z3/z1/z1/_1_  (.A(\v0/z2/z3/z1/temp [1]),
    .B(\v0/z2/z3/z1/temp [0]),
    .X(\v0/z2/q2 [1]));
 sky130_fd_sc_hd__and2_0 \v0/z2/z3/z1/z2/_0_  (.A(\v0/z2/z3/z1/temp [3]),
    .B(\v0/z2/z3/z1/temp [2]),
    .X(\v0/z2/z3/q0 [3]));
 sky130_fd_sc_hd__xor2_1 \v0/z2/z3/z1/z2/_1_  (.A(\v0/z2/z3/z1/temp [3]),
    .B(\v0/z2/z3/z1/temp [2]),
    .X(\v0/z2/z3/q0 [2]));
 sky130_fd_sc_hd__and2_0 \v0/z2/z3/z2/_0_  (.A(abs_b[4]),
    .B(abs_a[10]),
    .X(\v0/z2/z3/q1 [0]));
 sky130_fd_sc_hd__and2_0 \v0/z2/z3/z2/_1_  (.A(abs_b[4]),
    .B(abs_a[11]),
    .X(\v0/z2/z3/z2/temp [0]));
 sky130_fd_sc_hd__and2_0 \v0/z2/z3/z2/_2_  (.A(abs_a[10]),
    .B(abs_b[5]),
    .X(\v0/z2/z3/z2/temp [1]));
 sky130_fd_sc_hd__and2_0 \v0/z2/z3/z2/_3_  (.A(abs_a[11]),
    .B(abs_b[5]),
    .X(\v0/z2/z3/z2/temp [2]));
 sky130_fd_sc_hd__and2_0 \v0/z2/z3/z2/z1/_0_  (.A(\v0/z2/z3/z2/temp [1]),
    .B(\v0/z2/z3/z2/temp [0]),
    .X(\v0/z2/z3/z2/temp [3]));
 sky130_fd_sc_hd__xor2_1 \v0/z2/z3/z2/z1/_1_  (.A(\v0/z2/z3/z2/temp [1]),
    .B(\v0/z2/z3/z2/temp [0]),
    .X(\v0/z2/z3/q1 [1]));
 sky130_fd_sc_hd__and2_0 \v0/z2/z3/z2/z2/_0_  (.A(\v0/z2/z3/z2/temp [3]),
    .B(\v0/z2/z3/z2/temp [2]),
    .X(\v0/z2/z3/q1 [3]));
 sky130_fd_sc_hd__xor2_1 \v0/z2/z3/z2/z2/_1_  (.A(\v0/z2/z3/z2/temp [3]),
    .B(\v0/z2/z3/z2/temp [2]),
    .X(\v0/z2/z3/q1 [2]));
 sky130_fd_sc_hd__and2_0 \v0/z2/z3/z3/_0_  (.A(abs_b[6]),
    .B(abs_a[8]),
    .X(\v0/z2/z3/q2 [0]));
 sky130_fd_sc_hd__and2_0 \v0/z2/z3/z3/_1_  (.A(abs_b[6]),
    .B(abs_a[9]),
    .X(\v0/z2/z3/z3/temp [0]));
 sky130_fd_sc_hd__and2_0 \v0/z2/z3/z3/_2_  (.A(abs_a[8]),
    .B(abs_b[7]),
    .X(\v0/z2/z3/z3/temp [1]));
 sky130_fd_sc_hd__and2_0 \v0/z2/z3/z3/_3_  (.A(abs_a[9]),
    .B(abs_b[7]),
    .X(\v0/z2/z3/z3/temp [2]));
 sky130_fd_sc_hd__and2_0 \v0/z2/z3/z3/z1/_0_  (.A(\v0/z2/z3/z3/temp [1]),
    .B(\v0/z2/z3/z3/temp [0]),
    .X(\v0/z2/z3/z3/temp [3]));
 sky130_fd_sc_hd__xor2_1 \v0/z2/z3/z3/z1/_1_  (.A(\v0/z2/z3/z3/temp [1]),
    .B(\v0/z2/z3/z3/temp [0]),
    .X(\v0/z2/z3/q2 [1]));
 sky130_fd_sc_hd__and2_0 \v0/z2/z3/z3/z2/_0_  (.A(\v0/z2/z3/z3/temp [3]),
    .B(\v0/z2/z3/z3/temp [2]),
    .X(\v0/z2/z3/q2 [3]));
 sky130_fd_sc_hd__xor2_1 \v0/z2/z3/z3/z2/_1_  (.A(\v0/z2/z3/z3/temp [3]),
    .B(\v0/z2/z3/z3/temp [2]),
    .X(\v0/z2/z3/q2 [2]));
 sky130_fd_sc_hd__and2_0 \v0/z2/z3/z4/_0_  (.A(abs_b[6]),
    .B(abs_a[10]),
    .X(\v0/z2/z3/q3 [0]));
 sky130_fd_sc_hd__and2_0 \v0/z2/z3/z4/_1_  (.A(abs_b[6]),
    .B(abs_a[11]),
    .X(\v0/z2/z3/z4/temp [0]));
 sky130_fd_sc_hd__and2_0 \v0/z2/z3/z4/_2_  (.A(abs_a[10]),
    .B(abs_b[7]),
    .X(\v0/z2/z3/z4/temp [1]));
 sky130_fd_sc_hd__and2_0 \v0/z2/z3/z4/_3_  (.A(abs_a[11]),
    .B(abs_b[7]),
    .X(\v0/z2/z3/z4/temp [2]));
 sky130_fd_sc_hd__and2_0 \v0/z2/z3/z4/z1/_0_  (.A(\v0/z2/z3/z4/temp [1]),
    .B(\v0/z2/z3/z4/temp [0]),
    .X(\v0/z2/z3/z4/temp [3]));
 sky130_fd_sc_hd__xor2_1 \v0/z2/z3/z4/z1/_1_  (.A(\v0/z2/z3/z4/temp [1]),
    .B(\v0/z2/z3/z4/temp [0]),
    .X(\v0/z2/z3/q3 [1]));
 sky130_fd_sc_hd__and2_0 \v0/z2/z3/z4/z2/_0_  (.A(\v0/z2/z3/z4/temp [3]),
    .B(\v0/z2/z3/z4/temp [2]),
    .X(\v0/z2/z3/q3 [3]));
 sky130_fd_sc_hd__xor2_1 \v0/z2/z3/z4/z2/_1_  (.A(\v0/z2/z3/z4/temp [3]),
    .B(\v0/z2/z3/z4/temp [2]),
    .X(\v0/z2/z3/q3 [2]));
 sky130_fd_sc_hd__xnor2_1 \v0/z2/z3/z5/_07_  (.A(\v0/z2/z3/q0 [2]),
    .B(\v0/z2/z3/q1 [0]),
    .Y(\v0/z2/z3/z5/_00_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z2/z3/z5/_08_  (.A(\v0/z2/z3/_02_ ),
    .B(\v0/z2/z3/z5/_00_ ),
    .Y(\v0/z2/z3/q4 [0]));
 sky130_fd_sc_hd__maj3_1 \v0/z2/z3/z5/_09_  (.A(\v0/z2/z3/q0 [2]),
    .B(\v0/z2/z3/q1 [0]),
    .C(\v0/z2/z3/_02_ ),
    .X(\v0/z2/z3/z5/_01_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z2/z3/z5/_10_  (.A(\v0/z2/z3/q0 [3]),
    .B(\v0/z2/z3/q1 [1]),
    .Y(\v0/z2/z3/z5/_02_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z2/z3/z5/_11_  (.A(\v0/z2/z3/z5/_01_ ),
    .B(\v0/z2/z3/z5/_02_ ),
    .Y(\v0/z2/z3/q4 [1]));
 sky130_fd_sc_hd__maj3_1 \v0/z2/z3/z5/_12_  (.A(\v0/z2/z3/q0 [3]),
    .B(\v0/z2/z3/q1 [1]),
    .C(\v0/z2/z3/z5/_01_ ),
    .X(\v0/z2/z3/z5/_03_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z2/z3/z5/_13_  (.A(\v0/z2/z3/_00_ ),
    .B(\v0/z2/z3/q1 [2]),
    .Y(\v0/z2/z3/z5/_04_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z2/z3/z5/_14_  (.A(\v0/z2/z3/z5/_03_ ),
    .B(\v0/z2/z3/z5/_04_ ),
    .Y(\v0/z2/z3/q4 [2]));
 sky130_fd_sc_hd__maj3_1 \v0/z2/z3/z5/_15_  (.A(\v0/z2/z3/_00_ ),
    .B(\v0/z2/z3/q1 [2]),
    .C(\v0/z2/z3/z5/_03_ ),
    .X(\v0/z2/z3/z5/_05_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z2/z3/z5/_16_  (.A(\v0/z2/z3/_01_ ),
    .B(\v0/z2/z3/q1 [3]),
    .Y(\v0/z2/z3/z5/_06_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z2/z3/z5/_17_  (.A(\v0/z2/z3/z5/_05_ ),
    .B(\v0/z2/z3/z5/_06_ ),
    .Y(\v0/z2/z3/q4 [3]));
 sky130_fd_sc_hd__maj3_1 \v0/z2/z3/z5/_18_  (.A(\v0/z2/z3/_01_ ),
    .B(\v0/z2/z3/q1 [3]),
    .C(\v0/z2/z3/z5/_05_ ),
    .X(\v0/z2/z3/z5/Cout ));
 sky130_fd_sc_hd__xnor2_1 \v0/z2/z3/z6/_19_  (.A(\v0/z2/z3/_05_ ),
    .B(\v0/z2/z3/q2 [0]),
    .Y(\v0/z2/z3/z6/_00_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z2/z3/z6/_20_  (.A(\v0/z2/z3/_07_ ),
    .B(\v0/z2/z3/z6/_00_ ),
    .Y(\v0/z2/z3/q5 [0]));
 sky130_fd_sc_hd__maj3_1 \v0/z2/z3/z6/_21_  (.A(\v0/z2/z3/_05_ ),
    .B(\v0/z2/z3/q2 [0]),
    .C(\v0/z2/z3/_07_ ),
    .X(\v0/z2/z3/z6/_01_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z2/z3/z6/_22_  (.A(\v0/z2/z3/_06_ ),
    .B(\v0/z2/z3/q2 [1]),
    .Y(\v0/z2/z3/z6/_02_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z2/z3/z6/_23_  (.A(\v0/z2/z3/z6/_01_ ),
    .B(\v0/z2/z3/z6/_02_ ),
    .Y(\v0/z2/z3/q5 [1]));
 sky130_fd_sc_hd__maj3_1 \v0/z2/z3/z6/_24_  (.A(\v0/z2/z3/_06_ ),
    .B(\v0/z2/z3/q2 [1]),
    .C(\v0/z2/z3/z6/_01_ ),
    .X(\v0/z2/z3/z6/_03_ ));
 sky130_fd_sc_hd__lpflow_inputiso1p_1 \v0/z2/z3/z6/_25_  (.A(\v0/z2/z3/q3 [0]),
    .SLEEP(\v0/z2/z3/q2 [2]),
    .X(\v0/z2/z3/z6/_04_ ));
 sky130_fd_sc_hd__and2_0 \v0/z2/z3/z6/_26_  (.A(\v0/z2/z3/q3 [0]),
    .B(\v0/z2/z3/q2 [2]),
    .X(\v0/z2/z3/z6/_05_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z2/z3/z6/_27_  (.A(\v0/z2/z3/q3 [0]),
    .B(\v0/z2/z3/q2 [2]),
    .Y(\v0/z2/z3/z6/_06_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z2/z3/z6/_28_  (.A(\v0/z2/z3/z6/_04_ ),
    .B(\v0/z2/z3/z6/_06_ ),
    .Y(\v0/z2/z3/z6/_07_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z2/z3/z6/_29_  (.A(\v0/z2/z3/z6/_03_ ),
    .B(\v0/z2/z3/z6/_07_ ),
    .Y(\v0/z2/z3/q5 [2]));
 sky130_fd_sc_hd__nand2_1 \v0/z2/z3/z6/_30_  (.A(\v0/z2/z3/q3 [1]),
    .B(\v0/z2/z3/q2 [3]),
    .Y(\v0/z2/z3/z6/_08_ ));
 sky130_fd_sc_hd__xor2_1 \v0/z2/z3/z6/_31_  (.A(\v0/z2/z3/q3 [1]),
    .B(\v0/z2/z3/q2 [3]),
    .X(\v0/z2/z3/z6/_09_ ));
 sky130_fd_sc_hd__o21ai_0 \v0/z2/z3/z6/_32_  (.A1(\v0/z2/z3/z6/_03_ ),
    .A2(\v0/z2/z3/z6/_05_ ),
    .B1(\v0/z2/z3/z6/_04_ ),
    .Y(\v0/z2/z3/z6/_10_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z2/z3/z6/_33_  (.A(\v0/z2/z3/z6/_09_ ),
    .B(\v0/z2/z3/z6/_10_ ),
    .Y(\v0/z2/z3/q5 [3]));
 sky130_fd_sc_hd__nor2_1 \v0/z2/z3/z6/_34_  (.A(\v0/z2/z3/q3 [2]),
    .B(\v0/z2/z3/_03_ ),
    .Y(\v0/z2/z3/z6/_11_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z2/z3/z6/_35_  (.A(\v0/z2/z3/q3 [2]),
    .B(\v0/z2/z3/_03_ ),
    .Y(\v0/z2/z3/z6/_12_ ));
 sky130_fd_sc_hd__nand2b_1 \v0/z2/z3/z6/_36_  (.A_N(\v0/z2/z3/z6/_11_ ),
    .B(\v0/z2/z3/z6/_12_ ),
    .Y(\v0/z2/z3/z6/_13_ ));
 sky130_fd_sc_hd__o221ai_1 \v0/z2/z3/z6/_37_  (.A1(\v0/z2/z3/q3 [1]),
    .A2(\v0/z2/z3/q2 [3]),
    .B1(\v0/z2/z3/z6/_03_ ),
    .B2(\v0/z2/z3/z6/_05_ ),
    .C1(\v0/z2/z3/z6/_04_ ),
    .Y(\v0/z2/z3/z6/_14_ ));
 sky130_fd_sc_hd__a21oi_1 \v0/z2/z3/z6/_38_  (.A1(\v0/z2/z3/z6/_08_ ),
    .A2(\v0/z2/z3/z6/_14_ ),
    .B1(\v0/z2/z3/z6/_13_ ),
    .Y(\v0/z2/z3/z6/_15_ ));
 sky130_fd_sc_hd__and3_1 \v0/z2/z3/z6/_39_  (.A(\v0/z2/z3/z6/_08_ ),
    .B(\v0/z2/z3/z6/_13_ ),
    .C(\v0/z2/z3/z6/_14_ ),
    .X(\v0/z2/z3/z6/_16_ ));
 sky130_fd_sc_hd__nor2_1 \v0/z2/z3/z6/_40_  (.A(\v0/z2/z3/z6/_15_ ),
    .B(\v0/z2/z3/z6/_16_ ),
    .Y(\v0/z2/z3/q5 [4]));
 sky130_fd_sc_hd__xnor2_1 \v0/z2/z3/z6/_41_  (.A(\v0/z2/z3/q3 [3]),
    .B(\v0/z2/z3/_04_ ),
    .Y(\v0/z2/z3/z6/_17_ ));
 sky130_fd_sc_hd__a31oi_1 \v0/z2/z3/z6/_42_  (.A1(\v0/z2/z3/z6/_08_ ),
    .A2(\v0/z2/z3/z6/_12_ ),
    .A3(\v0/z2/z3/z6/_14_ ),
    .B1(\v0/z2/z3/z6/_11_ ),
    .Y(\v0/z2/z3/z6/_18_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z2/z3/z6/_43_  (.A(\v0/z2/z3/z6/_17_ ),
    .B(\v0/z2/z3/z6/_18_ ),
    .Y(\v0/z2/z3/q5 [5]));
 sky130_fd_sc_hd__maj3_1 \v0/z2/z3/z6/_44_  (.A(\v0/z2/z3/q3 [3]),
    .B(\v0/z2/z3/_04_ ),
    .C(\v0/z2/z3/z6/_18_ ),
    .X(\v0/z2/z3/z6/Cout ));
 sky130_fd_sc_hd__xnor2_1 \v0/z2/z3/z7/_19_  (.A(\v0/z2/z3/q5 [0]),
    .B(\v0/z2/z3/q4 [0]),
    .Y(\v0/z2/z3/z7/_00_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z2/z3/z7/_20_  (.A(\v0/z2/z3/_10_ ),
    .B(\v0/z2/z3/z7/_00_ ),
    .Y(\v0/z2/q2 [2]));
 sky130_fd_sc_hd__maj3_1 \v0/z2/z3/z7/_21_  (.A(\v0/z2/z3/q5 [0]),
    .B(\v0/z2/z3/q4 [0]),
    .C(\v0/z2/z3/_10_ ),
    .X(\v0/z2/z3/z7/_01_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z2/z3/z7/_22_  (.A(\v0/z2/z3/q5 [1]),
    .B(\v0/z2/z3/q4 [1]),
    .Y(\v0/z2/z3/z7/_02_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z2/z3/z7/_23_  (.A(\v0/z2/z3/z7/_01_ ),
    .B(\v0/z2/z3/z7/_02_ ),
    .Y(\v0/z2/q2 [3]));
 sky130_fd_sc_hd__maj3_1 \v0/z2/z3/z7/_24_  (.A(\v0/z2/z3/q5 [1]),
    .B(\v0/z2/z3/q4 [1]),
    .C(\v0/z2/z3/z7/_01_ ),
    .X(\v0/z2/z3/z7/_03_ ));
 sky130_fd_sc_hd__lpflow_inputiso1p_1 \v0/z2/z3/z7/_25_  (.A(\v0/z2/z3/q5 [2]),
    .SLEEP(\v0/z2/z3/q4 [2]),
    .X(\v0/z2/z3/z7/_04_ ));
 sky130_fd_sc_hd__and2_0 \v0/z2/z3/z7/_26_  (.A(\v0/z2/z3/q5 [2]),
    .B(\v0/z2/z3/q4 [2]),
    .X(\v0/z2/z3/z7/_05_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z2/z3/z7/_27_  (.A(\v0/z2/z3/q5 [2]),
    .B(\v0/z2/z3/q4 [2]),
    .Y(\v0/z2/z3/z7/_06_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z2/z3/z7/_28_  (.A(\v0/z2/z3/z7/_04_ ),
    .B(\v0/z2/z3/z7/_06_ ),
    .Y(\v0/z2/z3/z7/_07_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z2/z3/z7/_29_  (.A(\v0/z2/z3/z7/_03_ ),
    .B(\v0/z2/z3/z7/_07_ ),
    .Y(\v0/z2/q2 [4]));
 sky130_fd_sc_hd__nand2_1 \v0/z2/z3/z7/_30_  (.A(\v0/z2/z3/q5 [3]),
    .B(\v0/z2/z3/q4 [3]),
    .Y(\v0/z2/z3/z7/_08_ ));
 sky130_fd_sc_hd__xor2_1 \v0/z2/z3/z7/_31_  (.A(\v0/z2/z3/q5 [3]),
    .B(\v0/z2/z3/q4 [3]),
    .X(\v0/z2/z3/z7/_09_ ));
 sky130_fd_sc_hd__o21ai_0 \v0/z2/z3/z7/_32_  (.A1(\v0/z2/z3/z7/_03_ ),
    .A2(\v0/z2/z3/z7/_05_ ),
    .B1(\v0/z2/z3/z7/_04_ ),
    .Y(\v0/z2/z3/z7/_10_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z2/z3/z7/_33_  (.A(\v0/z2/z3/z7/_09_ ),
    .B(\v0/z2/z3/z7/_10_ ),
    .Y(\v0/z2/q2 [5]));
 sky130_fd_sc_hd__nor2_1 \v0/z2/z3/z7/_34_  (.A(\v0/z2/z3/q5 [4]),
    .B(\v0/z2/z3/_08_ ),
    .Y(\v0/z2/z3/z7/_11_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z2/z3/z7/_35_  (.A(\v0/z2/z3/q5 [4]),
    .B(\v0/z2/z3/_08_ ),
    .Y(\v0/z2/z3/z7/_12_ ));
 sky130_fd_sc_hd__nand2b_1 \v0/z2/z3/z7/_36_  (.A_N(\v0/z2/z3/z7/_11_ ),
    .B(\v0/z2/z3/z7/_12_ ),
    .Y(\v0/z2/z3/z7/_13_ ));
 sky130_fd_sc_hd__o221ai_1 \v0/z2/z3/z7/_37_  (.A1(\v0/z2/z3/q5 [3]),
    .A2(\v0/z2/z3/q4 [3]),
    .B1(\v0/z2/z3/z7/_03_ ),
    .B2(\v0/z2/z3/z7/_05_ ),
    .C1(\v0/z2/z3/z7/_04_ ),
    .Y(\v0/z2/z3/z7/_14_ ));
 sky130_fd_sc_hd__a21oi_1 \v0/z2/z3/z7/_38_  (.A1(\v0/z2/z3/z7/_08_ ),
    .A2(\v0/z2/z3/z7/_14_ ),
    .B1(\v0/z2/z3/z7/_13_ ),
    .Y(\v0/z2/z3/z7/_15_ ));
 sky130_fd_sc_hd__and3_1 \v0/z2/z3/z7/_39_  (.A(\v0/z2/z3/z7/_08_ ),
    .B(\v0/z2/z3/z7/_13_ ),
    .C(\v0/z2/z3/z7/_14_ ),
    .X(\v0/z2/z3/z7/_16_ ));
 sky130_fd_sc_hd__nor2_1 \v0/z2/z3/z7/_40_  (.A(\v0/z2/z3/z7/_15_ ),
    .B(\v0/z2/z3/z7/_16_ ),
    .Y(\v0/z2/q2 [6]));
 sky130_fd_sc_hd__xnor2_1 \v0/z2/z3/z7/_41_  (.A(\v0/z2/z3/q5 [5]),
    .B(\v0/z2/z3/_09_ ),
    .Y(\v0/z2/z3/z7/_17_ ));
 sky130_fd_sc_hd__a31oi_1 \v0/z2/z3/z7/_42_  (.A1(\v0/z2/z3/z7/_08_ ),
    .A2(\v0/z2/z3/z7/_12_ ),
    .A3(\v0/z2/z3/z7/_14_ ),
    .B1(\v0/z2/z3/z7/_11_ ),
    .Y(\v0/z2/z3/z7/_18_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z2/z3/z7/_43_  (.A(\v0/z2/z3/z7/_17_ ),
    .B(\v0/z2/z3/z7/_18_ ),
    .Y(\v0/z2/q2 [7]));
 sky130_fd_sc_hd__maj3_1 \v0/z2/z3/z7/_44_  (.A(\v0/z2/z3/q5 [5]),
    .B(\v0/z2/z3/_09_ ),
    .C(\v0/z2/z3/z7/_18_ ),
    .X(\v0/z2/z3/z7/Cout ));
 sky130_fd_sc_hd__conb_1 \v0/z2/z4/_11_  (.LO(\v0/z2/z4/_00_ ));
 sky130_fd_sc_hd__conb_1 \v0/z2/z4/_12_  (.LO(\v0/z2/z4/_01_ ));
 sky130_fd_sc_hd__conb_1 \v0/z2/z4/_13_  (.LO(\v0/z2/z4/_02_ ));
 sky130_fd_sc_hd__conb_1 \v0/z2/z4/_14_  (.LO(\v0/z2/z4/_03_ ));
 sky130_fd_sc_hd__conb_1 \v0/z2/z4/_15_  (.LO(\v0/z2/z4/_04_ ));
 sky130_fd_sc_hd__conb_1 \v0/z2/z4/_16_  (.LO(\v0/z2/z4/_05_ ));
 sky130_fd_sc_hd__conb_1 \v0/z2/z4/_17_  (.LO(\v0/z2/z4/_06_ ));
 sky130_fd_sc_hd__conb_1 \v0/z2/z4/_18_  (.LO(\v0/z2/z4/_07_ ));
 sky130_fd_sc_hd__conb_1 \v0/z2/z4/_19_  (.LO(\v0/z2/z4/_08_ ));
 sky130_fd_sc_hd__conb_1 \v0/z2/z4/_20_  (.LO(\v0/z2/z4/_09_ ));
 sky130_fd_sc_hd__conb_1 \v0/z2/z4/_21_  (.LO(\v0/z2/z4/_10_ ));
 sky130_fd_sc_hd__and2_0 \v0/z2/z4/z1/_0_  (.A(abs_b[4]),
    .B(abs_a[12]),
    .X(\v0/z2/q3 [0]));
 sky130_fd_sc_hd__and2_0 \v0/z2/z4/z1/_1_  (.A(abs_b[4]),
    .B(abs_a[13]),
    .X(\v0/z2/z4/z1/temp [0]));
 sky130_fd_sc_hd__and2_0 \v0/z2/z4/z1/_2_  (.A(abs_a[12]),
    .B(abs_b[5]),
    .X(\v0/z2/z4/z1/temp [1]));
 sky130_fd_sc_hd__and2_0 \v0/z2/z4/z1/_3_  (.A(abs_a[13]),
    .B(abs_b[5]),
    .X(\v0/z2/z4/z1/temp [2]));
 sky130_fd_sc_hd__and2_0 \v0/z2/z4/z1/z1/_0_  (.A(\v0/z2/z4/z1/temp [1]),
    .B(\v0/z2/z4/z1/temp [0]),
    .X(\v0/z2/z4/z1/temp [3]));
 sky130_fd_sc_hd__xor2_1 \v0/z2/z4/z1/z1/_1_  (.A(\v0/z2/z4/z1/temp [1]),
    .B(\v0/z2/z4/z1/temp [0]),
    .X(\v0/z2/q3 [1]));
 sky130_fd_sc_hd__and2_0 \v0/z2/z4/z1/z2/_0_  (.A(\v0/z2/z4/z1/temp [3]),
    .B(\v0/z2/z4/z1/temp [2]),
    .X(\v0/z2/z4/q0 [3]));
 sky130_fd_sc_hd__xor2_1 \v0/z2/z4/z1/z2/_1_  (.A(\v0/z2/z4/z1/temp [3]),
    .B(\v0/z2/z4/z1/temp [2]),
    .X(\v0/z2/z4/q0 [2]));
 sky130_fd_sc_hd__and2_0 \v0/z2/z4/z2/_0_  (.A(abs_b[4]),
    .B(abs_a[14]),
    .X(\v0/z2/z4/q1 [0]));
 sky130_fd_sc_hd__and2_0 \v0/z2/z4/z2/_1_  (.A(abs_b[4]),
    .B(abs_a[15]),
    .X(\v0/z2/z4/z2/temp [0]));
 sky130_fd_sc_hd__and2_0 \v0/z2/z4/z2/_2_  (.A(abs_a[14]),
    .B(abs_b[5]),
    .X(\v0/z2/z4/z2/temp [1]));
 sky130_fd_sc_hd__and2_0 \v0/z2/z4/z2/_3_  (.A(abs_a[15]),
    .B(abs_b[5]),
    .X(\v0/z2/z4/z2/temp [2]));
 sky130_fd_sc_hd__and2_0 \v0/z2/z4/z2/z1/_0_  (.A(\v0/z2/z4/z2/temp [1]),
    .B(\v0/z2/z4/z2/temp [0]),
    .X(\v0/z2/z4/z2/temp [3]));
 sky130_fd_sc_hd__xor2_1 \v0/z2/z4/z2/z1/_1_  (.A(\v0/z2/z4/z2/temp [1]),
    .B(\v0/z2/z4/z2/temp [0]),
    .X(\v0/z2/z4/q1 [1]));
 sky130_fd_sc_hd__and2_0 \v0/z2/z4/z2/z2/_0_  (.A(\v0/z2/z4/z2/temp [3]),
    .B(\v0/z2/z4/z2/temp [2]),
    .X(\v0/z2/z4/q1 [3]));
 sky130_fd_sc_hd__xor2_1 \v0/z2/z4/z2/z2/_1_  (.A(\v0/z2/z4/z2/temp [3]),
    .B(\v0/z2/z4/z2/temp [2]),
    .X(\v0/z2/z4/q1 [2]));
 sky130_fd_sc_hd__and2_0 \v0/z2/z4/z3/_0_  (.A(abs_b[6]),
    .B(abs_a[12]),
    .X(\v0/z2/z4/q2 [0]));
 sky130_fd_sc_hd__and2_0 \v0/z2/z4/z3/_1_  (.A(abs_b[6]),
    .B(abs_a[13]),
    .X(\v0/z2/z4/z3/temp [0]));
 sky130_fd_sc_hd__and2_0 \v0/z2/z4/z3/_2_  (.A(abs_a[12]),
    .B(abs_b[7]),
    .X(\v0/z2/z4/z3/temp [1]));
 sky130_fd_sc_hd__and2_0 \v0/z2/z4/z3/_3_  (.A(abs_a[13]),
    .B(abs_b[7]),
    .X(\v0/z2/z4/z3/temp [2]));
 sky130_fd_sc_hd__and2_0 \v0/z2/z4/z3/z1/_0_  (.A(\v0/z2/z4/z3/temp [1]),
    .B(\v0/z2/z4/z3/temp [0]),
    .X(\v0/z2/z4/z3/temp [3]));
 sky130_fd_sc_hd__xor2_1 \v0/z2/z4/z3/z1/_1_  (.A(\v0/z2/z4/z3/temp [1]),
    .B(\v0/z2/z4/z3/temp [0]),
    .X(\v0/z2/z4/q2 [1]));
 sky130_fd_sc_hd__and2_0 \v0/z2/z4/z3/z2/_0_  (.A(\v0/z2/z4/z3/temp [3]),
    .B(\v0/z2/z4/z3/temp [2]),
    .X(\v0/z2/z4/q2 [3]));
 sky130_fd_sc_hd__xor2_1 \v0/z2/z4/z3/z2/_1_  (.A(\v0/z2/z4/z3/temp [3]),
    .B(\v0/z2/z4/z3/temp [2]),
    .X(\v0/z2/z4/q2 [2]));
 sky130_fd_sc_hd__and2_0 \v0/z2/z4/z4/_0_  (.A(abs_b[6]),
    .B(abs_a[14]),
    .X(\v0/z2/z4/q3 [0]));
 sky130_fd_sc_hd__and2_0 \v0/z2/z4/z4/_1_  (.A(abs_b[6]),
    .B(abs_a[15]),
    .X(\v0/z2/z4/z4/temp [0]));
 sky130_fd_sc_hd__and2_0 \v0/z2/z4/z4/_2_  (.A(abs_a[14]),
    .B(abs_b[7]),
    .X(\v0/z2/z4/z4/temp [1]));
 sky130_fd_sc_hd__and2_0 \v0/z2/z4/z4/_3_  (.A(abs_a[15]),
    .B(abs_b[7]),
    .X(\v0/z2/z4/z4/temp [2]));
 sky130_fd_sc_hd__and2_0 \v0/z2/z4/z4/z1/_0_  (.A(\v0/z2/z4/z4/temp [1]),
    .B(\v0/z2/z4/z4/temp [0]),
    .X(\v0/z2/z4/z4/temp [3]));
 sky130_fd_sc_hd__xor2_1 \v0/z2/z4/z4/z1/_1_  (.A(\v0/z2/z4/z4/temp [1]),
    .B(\v0/z2/z4/z4/temp [0]),
    .X(\v0/z2/z4/q3 [1]));
 sky130_fd_sc_hd__and2_0 \v0/z2/z4/z4/z2/_0_  (.A(\v0/z2/z4/z4/temp [3]),
    .B(\v0/z2/z4/z4/temp [2]),
    .X(\v0/z2/z4/q3 [3]));
 sky130_fd_sc_hd__xor2_1 \v0/z2/z4/z4/z2/_1_  (.A(\v0/z2/z4/z4/temp [3]),
    .B(\v0/z2/z4/z4/temp [2]),
    .X(\v0/z2/z4/q3 [2]));
 sky130_fd_sc_hd__xnor2_1 \v0/z2/z4/z5/_07_  (.A(\v0/z2/z4/q0 [2]),
    .B(\v0/z2/z4/q1 [0]),
    .Y(\v0/z2/z4/z5/_00_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z2/z4/z5/_08_  (.A(\v0/z2/z4/_02_ ),
    .B(\v0/z2/z4/z5/_00_ ),
    .Y(\v0/z2/z4/q4 [0]));
 sky130_fd_sc_hd__maj3_1 \v0/z2/z4/z5/_09_  (.A(\v0/z2/z4/q0 [2]),
    .B(\v0/z2/z4/q1 [0]),
    .C(\v0/z2/z4/_02_ ),
    .X(\v0/z2/z4/z5/_01_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z2/z4/z5/_10_  (.A(\v0/z2/z4/q0 [3]),
    .B(\v0/z2/z4/q1 [1]),
    .Y(\v0/z2/z4/z5/_02_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z2/z4/z5/_11_  (.A(\v0/z2/z4/z5/_01_ ),
    .B(\v0/z2/z4/z5/_02_ ),
    .Y(\v0/z2/z4/q4 [1]));
 sky130_fd_sc_hd__maj3_1 \v0/z2/z4/z5/_12_  (.A(\v0/z2/z4/q0 [3]),
    .B(\v0/z2/z4/q1 [1]),
    .C(\v0/z2/z4/z5/_01_ ),
    .X(\v0/z2/z4/z5/_03_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z2/z4/z5/_13_  (.A(\v0/z2/z4/_00_ ),
    .B(\v0/z2/z4/q1 [2]),
    .Y(\v0/z2/z4/z5/_04_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z2/z4/z5/_14_  (.A(\v0/z2/z4/z5/_03_ ),
    .B(\v0/z2/z4/z5/_04_ ),
    .Y(\v0/z2/z4/q4 [2]));
 sky130_fd_sc_hd__maj3_1 \v0/z2/z4/z5/_15_  (.A(\v0/z2/z4/_00_ ),
    .B(\v0/z2/z4/q1 [2]),
    .C(\v0/z2/z4/z5/_03_ ),
    .X(\v0/z2/z4/z5/_05_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z2/z4/z5/_16_  (.A(\v0/z2/z4/_01_ ),
    .B(\v0/z2/z4/q1 [3]),
    .Y(\v0/z2/z4/z5/_06_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z2/z4/z5/_17_  (.A(\v0/z2/z4/z5/_05_ ),
    .B(\v0/z2/z4/z5/_06_ ),
    .Y(\v0/z2/z4/q4 [3]));
 sky130_fd_sc_hd__maj3_1 \v0/z2/z4/z5/_18_  (.A(\v0/z2/z4/_01_ ),
    .B(\v0/z2/z4/q1 [3]),
    .C(\v0/z2/z4/z5/_05_ ),
    .X(\v0/z2/z4/z5/Cout ));
 sky130_fd_sc_hd__xnor2_1 \v0/z2/z4/z6/_19_  (.A(\v0/z2/z4/_05_ ),
    .B(\v0/z2/z4/q2 [0]),
    .Y(\v0/z2/z4/z6/_00_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z2/z4/z6/_20_  (.A(\v0/z2/z4/_07_ ),
    .B(\v0/z2/z4/z6/_00_ ),
    .Y(\v0/z2/z4/q5 [0]));
 sky130_fd_sc_hd__maj3_1 \v0/z2/z4/z6/_21_  (.A(\v0/z2/z4/_05_ ),
    .B(\v0/z2/z4/q2 [0]),
    .C(\v0/z2/z4/_07_ ),
    .X(\v0/z2/z4/z6/_01_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z2/z4/z6/_22_  (.A(\v0/z2/z4/_06_ ),
    .B(\v0/z2/z4/q2 [1]),
    .Y(\v0/z2/z4/z6/_02_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z2/z4/z6/_23_  (.A(\v0/z2/z4/z6/_01_ ),
    .B(\v0/z2/z4/z6/_02_ ),
    .Y(\v0/z2/z4/q5 [1]));
 sky130_fd_sc_hd__maj3_1 \v0/z2/z4/z6/_24_  (.A(\v0/z2/z4/_06_ ),
    .B(\v0/z2/z4/q2 [1]),
    .C(\v0/z2/z4/z6/_01_ ),
    .X(\v0/z2/z4/z6/_03_ ));
 sky130_fd_sc_hd__lpflow_inputiso1p_1 \v0/z2/z4/z6/_25_  (.A(\v0/z2/z4/q3 [0]),
    .SLEEP(\v0/z2/z4/q2 [2]),
    .X(\v0/z2/z4/z6/_04_ ));
 sky130_fd_sc_hd__and2_0 \v0/z2/z4/z6/_26_  (.A(\v0/z2/z4/q3 [0]),
    .B(\v0/z2/z4/q2 [2]),
    .X(\v0/z2/z4/z6/_05_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z2/z4/z6/_27_  (.A(\v0/z2/z4/q3 [0]),
    .B(\v0/z2/z4/q2 [2]),
    .Y(\v0/z2/z4/z6/_06_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z2/z4/z6/_28_  (.A(\v0/z2/z4/z6/_04_ ),
    .B(\v0/z2/z4/z6/_06_ ),
    .Y(\v0/z2/z4/z6/_07_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z2/z4/z6/_29_  (.A(\v0/z2/z4/z6/_03_ ),
    .B(\v0/z2/z4/z6/_07_ ),
    .Y(\v0/z2/z4/q5 [2]));
 sky130_fd_sc_hd__nand2_1 \v0/z2/z4/z6/_30_  (.A(\v0/z2/z4/q3 [1]),
    .B(\v0/z2/z4/q2 [3]),
    .Y(\v0/z2/z4/z6/_08_ ));
 sky130_fd_sc_hd__xor2_1 \v0/z2/z4/z6/_31_  (.A(\v0/z2/z4/q3 [1]),
    .B(\v0/z2/z4/q2 [3]),
    .X(\v0/z2/z4/z6/_09_ ));
 sky130_fd_sc_hd__o21ai_0 \v0/z2/z4/z6/_32_  (.A1(\v0/z2/z4/z6/_03_ ),
    .A2(\v0/z2/z4/z6/_05_ ),
    .B1(\v0/z2/z4/z6/_04_ ),
    .Y(\v0/z2/z4/z6/_10_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z2/z4/z6/_33_  (.A(\v0/z2/z4/z6/_09_ ),
    .B(\v0/z2/z4/z6/_10_ ),
    .Y(\v0/z2/z4/q5 [3]));
 sky130_fd_sc_hd__nor2_1 \v0/z2/z4/z6/_34_  (.A(\v0/z2/z4/q3 [2]),
    .B(\v0/z2/z4/_03_ ),
    .Y(\v0/z2/z4/z6/_11_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z2/z4/z6/_35_  (.A(\v0/z2/z4/q3 [2]),
    .B(\v0/z2/z4/_03_ ),
    .Y(\v0/z2/z4/z6/_12_ ));
 sky130_fd_sc_hd__nand2b_1 \v0/z2/z4/z6/_36_  (.A_N(\v0/z2/z4/z6/_11_ ),
    .B(\v0/z2/z4/z6/_12_ ),
    .Y(\v0/z2/z4/z6/_13_ ));
 sky130_fd_sc_hd__o221ai_1 \v0/z2/z4/z6/_37_  (.A1(\v0/z2/z4/q3 [1]),
    .A2(\v0/z2/z4/q2 [3]),
    .B1(\v0/z2/z4/z6/_03_ ),
    .B2(\v0/z2/z4/z6/_05_ ),
    .C1(\v0/z2/z4/z6/_04_ ),
    .Y(\v0/z2/z4/z6/_14_ ));
 sky130_fd_sc_hd__a21oi_1 \v0/z2/z4/z6/_38_  (.A1(\v0/z2/z4/z6/_08_ ),
    .A2(\v0/z2/z4/z6/_14_ ),
    .B1(\v0/z2/z4/z6/_13_ ),
    .Y(\v0/z2/z4/z6/_15_ ));
 sky130_fd_sc_hd__and3_1 \v0/z2/z4/z6/_39_  (.A(\v0/z2/z4/z6/_08_ ),
    .B(\v0/z2/z4/z6/_13_ ),
    .C(\v0/z2/z4/z6/_14_ ),
    .X(\v0/z2/z4/z6/_16_ ));
 sky130_fd_sc_hd__nor2_1 \v0/z2/z4/z6/_40_  (.A(\v0/z2/z4/z6/_15_ ),
    .B(\v0/z2/z4/z6/_16_ ),
    .Y(\v0/z2/z4/q5 [4]));
 sky130_fd_sc_hd__xnor2_1 \v0/z2/z4/z6/_41_  (.A(\v0/z2/z4/q3 [3]),
    .B(\v0/z2/z4/_04_ ),
    .Y(\v0/z2/z4/z6/_17_ ));
 sky130_fd_sc_hd__a31oi_1 \v0/z2/z4/z6/_42_  (.A1(\v0/z2/z4/z6/_08_ ),
    .A2(\v0/z2/z4/z6/_12_ ),
    .A3(\v0/z2/z4/z6/_14_ ),
    .B1(\v0/z2/z4/z6/_11_ ),
    .Y(\v0/z2/z4/z6/_18_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z2/z4/z6/_43_  (.A(\v0/z2/z4/z6/_17_ ),
    .B(\v0/z2/z4/z6/_18_ ),
    .Y(\v0/z2/z4/q5 [5]));
 sky130_fd_sc_hd__maj3_1 \v0/z2/z4/z6/_44_  (.A(\v0/z2/z4/q3 [3]),
    .B(\v0/z2/z4/_04_ ),
    .C(\v0/z2/z4/z6/_18_ ),
    .X(\v0/z2/z4/z6/Cout ));
 sky130_fd_sc_hd__xnor2_1 \v0/z2/z4/z7/_19_  (.A(\v0/z2/z4/q5 [0]),
    .B(\v0/z2/z4/q4 [0]),
    .Y(\v0/z2/z4/z7/_00_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z2/z4/z7/_20_  (.A(\v0/z2/z4/_10_ ),
    .B(\v0/z2/z4/z7/_00_ ),
    .Y(\v0/z2/q3 [2]));
 sky130_fd_sc_hd__maj3_1 \v0/z2/z4/z7/_21_  (.A(\v0/z2/z4/q5 [0]),
    .B(\v0/z2/z4/q4 [0]),
    .C(\v0/z2/z4/_10_ ),
    .X(\v0/z2/z4/z7/_01_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z2/z4/z7/_22_  (.A(\v0/z2/z4/q5 [1]),
    .B(\v0/z2/z4/q4 [1]),
    .Y(\v0/z2/z4/z7/_02_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z2/z4/z7/_23_  (.A(\v0/z2/z4/z7/_01_ ),
    .B(\v0/z2/z4/z7/_02_ ),
    .Y(\v0/z2/q3 [3]));
 sky130_fd_sc_hd__maj3_1 \v0/z2/z4/z7/_24_  (.A(\v0/z2/z4/q5 [1]),
    .B(\v0/z2/z4/q4 [1]),
    .C(\v0/z2/z4/z7/_01_ ),
    .X(\v0/z2/z4/z7/_03_ ));
 sky130_fd_sc_hd__lpflow_inputiso1p_1 \v0/z2/z4/z7/_25_  (.A(\v0/z2/z4/q5 [2]),
    .SLEEP(\v0/z2/z4/q4 [2]),
    .X(\v0/z2/z4/z7/_04_ ));
 sky130_fd_sc_hd__and2_0 \v0/z2/z4/z7/_26_  (.A(\v0/z2/z4/q5 [2]),
    .B(\v0/z2/z4/q4 [2]),
    .X(\v0/z2/z4/z7/_05_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z2/z4/z7/_27_  (.A(\v0/z2/z4/q5 [2]),
    .B(\v0/z2/z4/q4 [2]),
    .Y(\v0/z2/z4/z7/_06_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z2/z4/z7/_28_  (.A(\v0/z2/z4/z7/_04_ ),
    .B(\v0/z2/z4/z7/_06_ ),
    .Y(\v0/z2/z4/z7/_07_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z2/z4/z7/_29_  (.A(\v0/z2/z4/z7/_03_ ),
    .B(\v0/z2/z4/z7/_07_ ),
    .Y(\v0/z2/q3 [4]));
 sky130_fd_sc_hd__nand2_1 \v0/z2/z4/z7/_30_  (.A(\v0/z2/z4/q5 [3]),
    .B(\v0/z2/z4/q4 [3]),
    .Y(\v0/z2/z4/z7/_08_ ));
 sky130_fd_sc_hd__xor2_1 \v0/z2/z4/z7/_31_  (.A(\v0/z2/z4/q5 [3]),
    .B(\v0/z2/z4/q4 [3]),
    .X(\v0/z2/z4/z7/_09_ ));
 sky130_fd_sc_hd__o21ai_0 \v0/z2/z4/z7/_32_  (.A1(\v0/z2/z4/z7/_03_ ),
    .A2(\v0/z2/z4/z7/_05_ ),
    .B1(\v0/z2/z4/z7/_04_ ),
    .Y(\v0/z2/z4/z7/_10_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z2/z4/z7/_33_  (.A(\v0/z2/z4/z7/_09_ ),
    .B(\v0/z2/z4/z7/_10_ ),
    .Y(\v0/z2/q3 [5]));
 sky130_fd_sc_hd__nor2_1 \v0/z2/z4/z7/_34_  (.A(\v0/z2/z4/q5 [4]),
    .B(\v0/z2/z4/_08_ ),
    .Y(\v0/z2/z4/z7/_11_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z2/z4/z7/_35_  (.A(\v0/z2/z4/q5 [4]),
    .B(\v0/z2/z4/_08_ ),
    .Y(\v0/z2/z4/z7/_12_ ));
 sky130_fd_sc_hd__nand2b_1 \v0/z2/z4/z7/_36_  (.A_N(\v0/z2/z4/z7/_11_ ),
    .B(\v0/z2/z4/z7/_12_ ),
    .Y(\v0/z2/z4/z7/_13_ ));
 sky130_fd_sc_hd__o221ai_1 \v0/z2/z4/z7/_37_  (.A1(\v0/z2/z4/q5 [3]),
    .A2(\v0/z2/z4/q4 [3]),
    .B1(\v0/z2/z4/z7/_03_ ),
    .B2(\v0/z2/z4/z7/_05_ ),
    .C1(\v0/z2/z4/z7/_04_ ),
    .Y(\v0/z2/z4/z7/_14_ ));
 sky130_fd_sc_hd__a21oi_1 \v0/z2/z4/z7/_38_  (.A1(\v0/z2/z4/z7/_08_ ),
    .A2(\v0/z2/z4/z7/_14_ ),
    .B1(\v0/z2/z4/z7/_13_ ),
    .Y(\v0/z2/z4/z7/_15_ ));
 sky130_fd_sc_hd__and3_1 \v0/z2/z4/z7/_39_  (.A(\v0/z2/z4/z7/_08_ ),
    .B(\v0/z2/z4/z7/_13_ ),
    .C(\v0/z2/z4/z7/_14_ ),
    .X(\v0/z2/z4/z7/_16_ ));
 sky130_fd_sc_hd__nor2_1 \v0/z2/z4/z7/_40_  (.A(\v0/z2/z4/z7/_15_ ),
    .B(\v0/z2/z4/z7/_16_ ),
    .Y(\v0/z2/q3 [6]));
 sky130_fd_sc_hd__xnor2_1 \v0/z2/z4/z7/_41_  (.A(\v0/z2/z4/q5 [5]),
    .B(\v0/z2/z4/_09_ ),
    .Y(\v0/z2/z4/z7/_17_ ));
 sky130_fd_sc_hd__a31oi_1 \v0/z2/z4/z7/_42_  (.A1(\v0/z2/z4/z7/_08_ ),
    .A2(\v0/z2/z4/z7/_12_ ),
    .A3(\v0/z2/z4/z7/_14_ ),
    .B1(\v0/z2/z4/z7/_11_ ),
    .Y(\v0/z2/z4/z7/_18_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z2/z4/z7/_43_  (.A(\v0/z2/z4/z7/_17_ ),
    .B(\v0/z2/z4/z7/_18_ ),
    .Y(\v0/z2/q3 [7]));
 sky130_fd_sc_hd__maj3_1 \v0/z2/z4/z7/_44_  (.A(\v0/z2/z4/q5 [5]),
    .B(\v0/z2/z4/_09_ ),
    .C(\v0/z2/z4/z7/_18_ ),
    .X(\v0/z2/z4/z7/Cout ));
 sky130_fd_sc_hd__xnor2_1 \v0/z2/z5/_27_  (.A(\v0/z2/q0 [4]),
    .B(\v0/z2/q1 [0]),
    .Y(\v0/z2/z5/_00_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z2/z5/_28_  (.A(\v0/z2/_04_ ),
    .B(\v0/z2/z5/_00_ ),
    .Y(\v0/z2/q4 [0]));
 sky130_fd_sc_hd__maj3_1 \v0/z2/z5/_29_  (.A(\v0/z2/q0 [4]),
    .B(\v0/z2/q1 [0]),
    .C(\v0/z2/_04_ ),
    .X(\v0/z2/z5/_01_ ));
 sky130_fd_sc_hd__lpflow_inputiso1p_1 \v0/z2/z5/_30_  (.A(\v0/z2/q0 [5]),
    .SLEEP(\v0/z2/q1 [1]),
    .X(\v0/z2/z5/_02_ ));
 sky130_fd_sc_hd__and2_0 \v0/z2/z5/_31_  (.A(\v0/z2/q0 [5]),
    .B(\v0/z2/q1 [1]),
    .X(\v0/z2/z5/_03_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z2/z5/_32_  (.A(\v0/z2/q0 [5]),
    .B(\v0/z2/q1 [1]),
    .Y(\v0/z2/z5/_04_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z2/z5/_33_  (.A(\v0/z2/z5/_02_ ),
    .B(\v0/z2/z5/_04_ ),
    .Y(\v0/z2/z5/_05_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z2/z5/_34_  (.A(\v0/z2/z5/_01_ ),
    .B(\v0/z2/z5/_05_ ),
    .Y(\v0/z2/q4 [1]));
 sky130_fd_sc_hd__nand2_1 \v0/z2/z5/_35_  (.A(\v0/z2/q0 [6]),
    .B(\v0/z2/q1 [2]),
    .Y(\v0/z2/z5/_06_ ));
 sky130_fd_sc_hd__xor2_1 \v0/z2/z5/_36_  (.A(\v0/z2/q0 [6]),
    .B(\v0/z2/q1 [2]),
    .X(\v0/z2/z5/_07_ ));
 sky130_fd_sc_hd__o21ai_0 \v0/z2/z5/_37_  (.A1(\v0/z2/z5/_01_ ),
    .A2(\v0/z2/z5/_03_ ),
    .B1(\v0/z2/z5/_02_ ),
    .Y(\v0/z2/z5/_08_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z2/z5/_38_  (.A(\v0/z2/z5/_07_ ),
    .B(\v0/z2/z5/_08_ ),
    .Y(\v0/z2/q4 [2]));
 sky130_fd_sc_hd__nor2_1 \v0/z2/z5/_39_  (.A(\v0/z2/q0 [7]),
    .B(\v0/z2/q1 [3]),
    .Y(\v0/z2/z5/_09_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z2/z5/_40_  (.A(\v0/z2/q0 [7]),
    .B(\v0/z2/q1 [3]),
    .Y(\v0/z2/z5/_10_ ));
 sky130_fd_sc_hd__nor2b_1 \v0/z2/z5/_41_  (.A(\v0/z2/z5/_09_ ),
    .B_N(\v0/z2/z5/_10_ ),
    .Y(\v0/z2/z5/_11_ ));
 sky130_fd_sc_hd__o221ai_1 \v0/z2/z5/_42_  (.A1(\v0/z2/q0 [6]),
    .A2(\v0/z2/q1 [2]),
    .B1(\v0/z2/z5/_01_ ),
    .B2(\v0/z2/z5/_03_ ),
    .C1(\v0/z2/z5/_02_ ),
    .Y(\v0/z2/z5/_12_ ));
 sky130_fd_sc_hd__and2_0 \v0/z2/z5/_43_  (.A(\v0/z2/z5/_06_ ),
    .B(\v0/z2/z5/_12_ ),
    .X(\v0/z2/z5/_13_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z2/z5/_44_  (.A(\v0/z2/z5/_11_ ),
    .B(\v0/z2/z5/_13_ ),
    .Y(\v0/z2/q4 [3]));
 sky130_fd_sc_hd__nor2_1 \v0/z2/z5/_45_  (.A(\v0/z2/_00_ ),
    .B(\v0/z2/q1 [4]),
    .Y(\v0/z2/z5/_14_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z2/z5/_46_  (.A(\v0/z2/_00_ ),
    .B(\v0/z2/q1 [4]),
    .Y(\v0/z2/z5/_15_ ));
 sky130_fd_sc_hd__nand2b_1 \v0/z2/z5/_47_  (.A_N(\v0/z2/z5/_14_ ),
    .B(\v0/z2/z5/_15_ ),
    .Y(\v0/z2/z5/_16_ ));
 sky130_fd_sc_hd__a21oi_1 \v0/z2/z5/_48_  (.A1(\v0/z2/z5/_10_ ),
    .A2(\v0/z2/z5/_13_ ),
    .B1(\v0/z2/z5/_09_ ),
    .Y(\v0/z2/z5/_17_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z2/z5/_49_  (.A(\v0/z2/z5/_16_ ),
    .B(\v0/z2/z5/_17_ ),
    .Y(\v0/z2/q4 [4]));
 sky130_fd_sc_hd__a311o_1 \v0/z2/z5/_50_  (.A1(\v0/z2/z5/_06_ ),
    .A2(\v0/z2/z5/_10_ ),
    .A3(\v0/z2/z5/_12_ ),
    .B1(\v0/z2/z5/_14_ ),
    .C1(\v0/z2/z5/_09_ ),
    .X(\v0/z2/z5/_18_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z2/z5/_51_  (.A(\v0/z2/z5/_15_ ),
    .B(\v0/z2/z5/_18_ ),
    .Y(\v0/z2/z5/_19_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z2/z5/_52_  (.A(\v0/z2/_01_ ),
    .B(\v0/z2/q1 [5]),
    .Y(\v0/z2/z5/_20_ ));
 sky130_fd_sc_hd__nor2_1 \v0/z2/z5/_53_  (.A(\v0/z2/_01_ ),
    .B(\v0/z2/q1 [5]),
    .Y(\v0/z2/z5/_21_ ));
 sky130_fd_sc_hd__a31oi_1 \v0/z2/z5/_54_  (.A1(\v0/z2/z5/_15_ ),
    .A2(\v0/z2/z5/_18_ ),
    .A3(\v0/z2/z5/_20_ ),
    .B1(\v0/z2/z5/_21_ ),
    .Y(\v0/z2/z5/_22_ ));
 sky130_fd_sc_hd__a21bo_1 \v0/z2/z5/_55_  (.A1(\v0/z2/z5/_20_ ),
    .A2(\v0/z2/z5/_22_ ),
    .B1_N(\v0/z2/z5/_19_ ),
    .X(\v0/z2/z5/_23_ ));
 sky130_fd_sc_hd__o21ai_0 \v0/z2/z5/_56_  (.A1(\v0/z2/z5/_21_ ),
    .A2(\v0/z2/z5/_22_ ),
    .B1(\v0/z2/z5/_23_ ),
    .Y(\v0/z2/q4 [5]));
 sky130_fd_sc_hd__xnor2_1 \v0/z2/z5/_57_  (.A(\v0/z2/_02_ ),
    .B(\v0/z2/q1 [6]),
    .Y(\v0/z2/z5/_24_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z2/z5/_58_  (.A(\v0/z2/z5/_22_ ),
    .B(\v0/z2/z5/_24_ ),
    .Y(\v0/z2/q4 [6]));
 sky130_fd_sc_hd__xnor2_1 \v0/z2/z5/_59_  (.A(\v0/z2/_03_ ),
    .B(\v0/z2/q1 [7]),
    .Y(\v0/z2/z5/_25_ ));
 sky130_fd_sc_hd__maj3_1 \v0/z2/z5/_60_  (.A(\v0/z2/_02_ ),
    .B(\v0/z2/q1 [6]),
    .C(\v0/z2/z5/_22_ ),
    .X(\v0/z2/z5/_26_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z2/z5/_61_  (.A(\v0/z2/z5/_25_ ),
    .B(\v0/z2/z5/_26_ ),
    .Y(\v0/z2/q4 [7]));
 sky130_fd_sc_hd__maj3_1 \v0/z2/z5/_62_  (.A(\v0/z2/_03_ ),
    .B(\v0/z2/q1 [7]),
    .C(\v0/z2/z5/_26_ ),
    .X(\v0/z2/z5/Cout ));
 sky130_fd_sc_hd__xnor2_1 \v0/z2/z6/_050_  (.A(\v0/z2/_09_ ),
    .B(\v0/z2/q2 [0]),
    .Y(\v0/z2/z6/_000_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z2/z6/_051_  (.A(\v0/z2/_13_ ),
    .B(\v0/z2/z6/_000_ ),
    .Y(\v0/z2/q5 [0]));
 sky130_fd_sc_hd__maj3_1 \v0/z2/z6/_052_  (.A(\v0/z2/_09_ ),
    .B(\v0/z2/q2 [0]),
    .C(\v0/z2/_13_ ),
    .X(\v0/z2/z6/_001_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z2/z6/_053_  (.A(\v0/z2/_10_ ),
    .B(\v0/z2/q2 [1]),
    .Y(\v0/z2/z6/_002_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z2/z6/_054_  (.A(\v0/z2/z6/_001_ ),
    .B(\v0/z2/z6/_002_ ),
    .Y(\v0/z2/q5 [1]));
 sky130_fd_sc_hd__maj3_1 \v0/z2/z6/_055_  (.A(\v0/z2/_10_ ),
    .B(\v0/z2/q2 [1]),
    .C(\v0/z2/z6/_001_ ),
    .X(\v0/z2/z6/_003_ ));
 sky130_fd_sc_hd__lpflow_inputiso1p_1 \v0/z2/z6/_056_  (.A(\v0/z2/_11_ ),
    .SLEEP(\v0/z2/q2 [2]),
    .X(\v0/z2/z6/_004_ ));
 sky130_fd_sc_hd__and2_0 \v0/z2/z6/_057_  (.A(\v0/z2/_11_ ),
    .B(\v0/z2/q2 [2]),
    .X(\v0/z2/z6/_005_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z2/z6/_058_  (.A(\v0/z2/_11_ ),
    .B(\v0/z2/q2 [2]),
    .Y(\v0/z2/z6/_006_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z2/z6/_059_  (.A(\v0/z2/z6/_004_ ),
    .B(\v0/z2/z6/_006_ ),
    .Y(\v0/z2/z6/_007_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z2/z6/_060_  (.A(\v0/z2/z6/_003_ ),
    .B(\v0/z2/z6/_007_ ),
    .Y(\v0/z2/q5 [2]));
 sky130_fd_sc_hd__nor2_1 \v0/z2/z6/_061_  (.A(\v0/z2/_12_ ),
    .B(\v0/z2/q2 [3]),
    .Y(\v0/z2/z6/_008_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z2/z6/_062_  (.A(\v0/z2/_12_ ),
    .B(\v0/z2/q2 [3]),
    .Y(\v0/z2/z6/_009_ ));
 sky130_fd_sc_hd__clkinv_1 \v0/z2/z6/_063_  (.A(\v0/z2/z6/_009_ ),
    .Y(\v0/z2/z6/_010_ ));
 sky130_fd_sc_hd__nor2_1 \v0/z2/z6/_064_  (.A(\v0/z2/z6/_008_ ),
    .B(\v0/z2/z6/_010_ ),
    .Y(\v0/z2/z6/_011_ ));
 sky130_fd_sc_hd__o21ai_0 \v0/z2/z6/_065_  (.A1(\v0/z2/z6/_003_ ),
    .A2(\v0/z2/z6/_005_ ),
    .B1(\v0/z2/z6/_004_ ),
    .Y(\v0/z2/z6/_012_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z2/z6/_066_  (.A(\v0/z2/z6/_011_ ),
    .B(\v0/z2/z6/_012_ ),
    .Y(\v0/z2/q5 [3]));
 sky130_fd_sc_hd__lpflow_inputiso1p_1 \v0/z2/z6/_067_  (.A(\v0/z2/q3 [0]),
    .SLEEP(\v0/z2/q2 [4]),
    .X(\v0/z2/z6/_013_ ));
 sky130_fd_sc_hd__and2_0 \v0/z2/z6/_068_  (.A(\v0/z2/q3 [0]),
    .B(\v0/z2/q2 [4]),
    .X(\v0/z2/z6/_014_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z2/z6/_069_  (.A(\v0/z2/q3 [0]),
    .B(\v0/z2/q2 [4]),
    .Y(\v0/z2/z6/_015_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z2/z6/_070_  (.A(\v0/z2/z6/_013_ ),
    .B(\v0/z2/z6/_015_ ),
    .Y(\v0/z2/z6/_016_ ));
 sky130_fd_sc_hd__o221a_1 \v0/z2/z6/_071_  (.A1(\v0/z2/_12_ ),
    .A2(\v0/z2/q2 [3]),
    .B1(\v0/z2/z6/_003_ ),
    .B2(\v0/z2/z6/_005_ ),
    .C1(\v0/z2/z6/_004_ ),
    .X(\v0/z2/z6/_017_ ));
 sky130_fd_sc_hd__a21oi_1 \v0/z2/z6/_072_  (.A1(\v0/z2/z6/_009_ ),
    .A2(\v0/z2/z6/_012_ ),
    .B1(\v0/z2/z6/_008_ ),
    .Y(\v0/z2/z6/_018_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z2/z6/_073_  (.A(\v0/z2/z6/_016_ ),
    .B(\v0/z2/z6/_018_ ),
    .Y(\v0/z2/q5 [4]));
 sky130_fd_sc_hd__lpflow_inputiso1p_1 \v0/z2/z6/_074_  (.A(\v0/z2/q3 [1]),
    .SLEEP(\v0/z2/q2 [5]),
    .X(\v0/z2/z6/_019_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z2/z6/_075_  (.A(\v0/z2/q3 [1]),
    .B(\v0/z2/q2 [5]),
    .Y(\v0/z2/z6/_020_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z2/z6/_076_  (.A(\v0/z2/z6/_019_ ),
    .B(\v0/z2/z6/_020_ ),
    .Y(\v0/z2/z6/_021_ ));
 sky130_fd_sc_hd__o21ai_0 \v0/z2/z6/_077_  (.A1(\v0/z2/z6/_014_ ),
    .A2(\v0/z2/z6/_018_ ),
    .B1(\v0/z2/z6/_013_ ),
    .Y(\v0/z2/z6/_022_ ));
 sky130_fd_sc_hd__xor2_1 \v0/z2/z6/_078_  (.A(\v0/z2/z6/_021_ ),
    .B(\v0/z2/z6/_022_ ),
    .X(\v0/z2/q5 [5]));
 sky130_fd_sc_hd__nor2_1 \v0/z2/z6/_079_  (.A(\v0/z2/q3 [2]),
    .B(\v0/z2/q2 [6]),
    .Y(\v0/z2/z6/_023_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z2/z6/_080_  (.A(\v0/z2/q3 [2]),
    .B(\v0/z2/q2 [6]),
    .Y(\v0/z2/z6/_024_ ));
 sky130_fd_sc_hd__nor2b_1 \v0/z2/z6/_081_  (.A(\v0/z2/z6/_023_ ),
    .B_N(\v0/z2/z6/_024_ ),
    .Y(\v0/z2/z6/_025_ ));
 sky130_fd_sc_hd__o311ai_0 \v0/z2/z6/_082_  (.A1(\v0/z2/z6/_010_ ),
    .A2(\v0/z2/z6/_014_ ),
    .A3(\v0/z2/z6/_017_ ),
    .B1(\v0/z2/z6/_019_ ),
    .C1(\v0/z2/z6/_013_ ),
    .Y(\v0/z2/z6/_026_ ));
 sky130_fd_sc_hd__and2_0 \v0/z2/z6/_083_  (.A(\v0/z2/z6/_020_ ),
    .B(\v0/z2/z6/_026_ ),
    .X(\v0/z2/z6/_027_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z2/z6/_084_  (.A(\v0/z2/z6/_025_ ),
    .B(\v0/z2/z6/_027_ ),
    .Y(\v0/z2/q5 [6]));
 sky130_fd_sc_hd__nor2_1 \v0/z2/z6/_085_  (.A(\v0/z2/q3 [3]),
    .B(\v0/z2/q2 [7]),
    .Y(\v0/z2/z6/_028_ ));
 sky130_fd_sc_hd__and2_0 \v0/z2/z6/_086_  (.A(\v0/z2/q3 [3]),
    .B(\v0/z2/q2 [7]),
    .X(\v0/z2/z6/_029_ ));
 sky130_fd_sc_hd__nor2_1 \v0/z2/z6/_087_  (.A(\v0/z2/z6/_028_ ),
    .B(\v0/z2/z6/_029_ ),
    .Y(\v0/z2/z6/_030_ ));
 sky130_fd_sc_hd__a21oi_1 \v0/z2/z6/_088_  (.A1(\v0/z2/z6/_024_ ),
    .A2(\v0/z2/z6/_027_ ),
    .B1(\v0/z2/z6/_023_ ),
    .Y(\v0/z2/z6/_031_ ));
 sky130_fd_sc_hd__xor2_1 \v0/z2/z6/_089_  (.A(\v0/z2/z6/_030_ ),
    .B(\v0/z2/z6/_031_ ),
    .X(\v0/z2/q5 [7]));
 sky130_fd_sc_hd__lpflow_inputiso1p_1 \v0/z2/z6/_090_  (.A(\v0/z2/q3 [4]),
    .SLEEP(\v0/z2/_05_ ),
    .X(\v0/z2/z6/_032_ ));
 sky130_fd_sc_hd__and2_0 \v0/z2/z6/_091_  (.A(\v0/z2/q3 [4]),
    .B(\v0/z2/_05_ ),
    .X(\v0/z2/z6/_033_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z2/z6/_092_  (.A(\v0/z2/q3 [4]),
    .B(\v0/z2/_05_ ),
    .Y(\v0/z2/z6/_034_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z2/z6/_093_  (.A(\v0/z2/z6/_032_ ),
    .B(\v0/z2/z6/_034_ ),
    .Y(\v0/z2/z6/_035_ ));
 sky130_fd_sc_hd__a311oi_1 \v0/z2/z6/_094_  (.A1(\v0/z2/z6/_020_ ),
    .A2(\v0/z2/z6/_024_ ),
    .A3(\v0/z2/z6/_026_ ),
    .B1(\v0/z2/z6/_028_ ),
    .C1(\v0/z2/z6/_023_ ),
    .Y(\v0/z2/z6/_036_ ));
 sky130_fd_sc_hd__lpflow_inputiso1p_1 \v0/z2/z6/_095_  (.A(\v0/z2/z6/_029_ ),
    .SLEEP(\v0/z2/z6/_036_ ),
    .X(\v0/z2/z6/_037_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z2/z6/_096_  (.A(\v0/z2/z6/_035_ ),
    .B(\v0/z2/z6/_037_ ),
    .Y(\v0/z2/q5 [8]));
 sky130_fd_sc_hd__lpflow_inputiso1p_1 \v0/z2/z6/_097_  (.A(\v0/z2/q3 [5]),
    .SLEEP(\v0/z2/_06_ ),
    .X(\v0/z2/z6/_038_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z2/z6/_098_  (.A(\v0/z2/q3 [5]),
    .B(\v0/z2/_06_ ),
    .Y(\v0/z2/z6/_039_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z2/z6/_099_  (.A(\v0/z2/z6/_038_ ),
    .B(\v0/z2/z6/_039_ ),
    .Y(\v0/z2/z6/_040_ ));
 sky130_fd_sc_hd__o21ai_0 \v0/z2/z6/_100_  (.A1(\v0/z2/z6/_033_ ),
    .A2(\v0/z2/z6/_037_ ),
    .B1(\v0/z2/z6/_032_ ),
    .Y(\v0/z2/z6/_041_ ));
 sky130_fd_sc_hd__xor2_1 \v0/z2/z6/_101_  (.A(\v0/z2/z6/_040_ ),
    .B(\v0/z2/z6/_041_ ),
    .X(\v0/z2/q5 [9]));
 sky130_fd_sc_hd__nor2_1 \v0/z2/z6/_102_  (.A(\v0/z2/q3 [6]),
    .B(\v0/z2/_07_ ),
    .Y(\v0/z2/z6/_042_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z2/z6/_103_  (.A(\v0/z2/q3 [6]),
    .B(\v0/z2/_07_ ),
    .Y(\v0/z2/z6/_043_ ));
 sky130_fd_sc_hd__nand2b_1 \v0/z2/z6/_104_  (.A_N(\v0/z2/z6/_042_ ),
    .B(\v0/z2/z6/_043_ ),
    .Y(\v0/z2/z6/_044_ ));
 sky130_fd_sc_hd__o311ai_0 \v0/z2/z6/_105_  (.A1(\v0/z2/z6/_029_ ),
    .A2(\v0/z2/z6/_033_ ),
    .A3(\v0/z2/z6/_036_ ),
    .B1(\v0/z2/z6/_038_ ),
    .C1(\v0/z2/z6/_032_ ),
    .Y(\v0/z2/z6/_045_ ));
 sky130_fd_sc_hd__a21oi_1 \v0/z2/z6/_106_  (.A1(\v0/z2/z6/_039_ ),
    .A2(\v0/z2/z6/_045_ ),
    .B1(\v0/z2/z6/_044_ ),
    .Y(\v0/z2/z6/_046_ ));
 sky130_fd_sc_hd__and3_1 \v0/z2/z6/_107_  (.A(\v0/z2/z6/_039_ ),
    .B(\v0/z2/z6/_044_ ),
    .C(\v0/z2/z6/_045_ ),
    .X(\v0/z2/z6/_047_ ));
 sky130_fd_sc_hd__nor2_1 \v0/z2/z6/_108_  (.A(\v0/z2/z6/_046_ ),
    .B(\v0/z2/z6/_047_ ),
    .Y(\v0/z2/q5 [10]));
 sky130_fd_sc_hd__xnor2_1 \v0/z2/z6/_109_  (.A(\v0/z2/q3 [7]),
    .B(\v0/z2/_08_ ),
    .Y(\v0/z2/z6/_048_ ));
 sky130_fd_sc_hd__a31oi_1 \v0/z2/z6/_110_  (.A1(\v0/z2/z6/_039_ ),
    .A2(\v0/z2/z6/_043_ ),
    .A3(\v0/z2/z6/_045_ ),
    .B1(\v0/z2/z6/_042_ ),
    .Y(\v0/z2/z6/_049_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z2/z6/_111_  (.A(\v0/z2/z6/_048_ ),
    .B(\v0/z2/z6/_049_ ),
    .Y(\v0/z2/q5 [11]));
 sky130_fd_sc_hd__maj3_1 \v0/z2/z6/_112_  (.A(\v0/z2/q3 [7]),
    .B(\v0/z2/_08_ ),
    .C(\v0/z2/z6/_049_ ),
    .X(\v0/z2/z6/Cout ));
 sky130_fd_sc_hd__xnor2_1 \v0/z2/z7/_050_  (.A(\v0/z2/q5 [0]),
    .B(\v0/z2/q4 [0]),
    .Y(\v0/z2/z7/_000_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z2/z7/_051_  (.A(\v0/z2/_18_ ),
    .B(\v0/z2/z7/_000_ ),
    .Y(\v0/q1 [4]));
 sky130_fd_sc_hd__maj3_1 \v0/z2/z7/_052_  (.A(\v0/z2/q5 [0]),
    .B(\v0/z2/q4 [0]),
    .C(\v0/z2/_18_ ),
    .X(\v0/z2/z7/_001_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z2/z7/_053_  (.A(\v0/z2/q5 [1]),
    .B(\v0/z2/q4 [1]),
    .Y(\v0/z2/z7/_002_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z2/z7/_054_  (.A(\v0/z2/z7/_001_ ),
    .B(\v0/z2/z7/_002_ ),
    .Y(\v0/q1 [5]));
 sky130_fd_sc_hd__maj3_1 \v0/z2/z7/_055_  (.A(\v0/z2/q5 [1]),
    .B(\v0/z2/q4 [1]),
    .C(\v0/z2/z7/_001_ ),
    .X(\v0/z2/z7/_003_ ));
 sky130_fd_sc_hd__lpflow_inputiso1p_1 \v0/z2/z7/_056_  (.A(\v0/z2/q5 [2]),
    .SLEEP(\v0/z2/q4 [2]),
    .X(\v0/z2/z7/_004_ ));
 sky130_fd_sc_hd__and2_0 \v0/z2/z7/_057_  (.A(\v0/z2/q5 [2]),
    .B(\v0/z2/q4 [2]),
    .X(\v0/z2/z7/_005_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z2/z7/_058_  (.A(\v0/z2/q5 [2]),
    .B(\v0/z2/q4 [2]),
    .Y(\v0/z2/z7/_006_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z2/z7/_059_  (.A(\v0/z2/z7/_004_ ),
    .B(\v0/z2/z7/_006_ ),
    .Y(\v0/z2/z7/_007_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z2/z7/_060_  (.A(\v0/z2/z7/_003_ ),
    .B(\v0/z2/z7/_007_ ),
    .Y(\v0/q1 [6]));
 sky130_fd_sc_hd__nor2_1 \v0/z2/z7/_061_  (.A(\v0/z2/q5 [3]),
    .B(\v0/z2/q4 [3]),
    .Y(\v0/z2/z7/_008_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z2/z7/_062_  (.A(\v0/z2/q5 [3]),
    .B(\v0/z2/q4 [3]),
    .Y(\v0/z2/z7/_009_ ));
 sky130_fd_sc_hd__clkinv_1 \v0/z2/z7/_063_  (.A(\v0/z2/z7/_009_ ),
    .Y(\v0/z2/z7/_010_ ));
 sky130_fd_sc_hd__nor2_1 \v0/z2/z7/_064_  (.A(\v0/z2/z7/_008_ ),
    .B(\v0/z2/z7/_010_ ),
    .Y(\v0/z2/z7/_011_ ));
 sky130_fd_sc_hd__o21ai_0 \v0/z2/z7/_065_  (.A1(\v0/z2/z7/_003_ ),
    .A2(\v0/z2/z7/_005_ ),
    .B1(\v0/z2/z7/_004_ ),
    .Y(\v0/z2/z7/_012_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z2/z7/_066_  (.A(\v0/z2/z7/_011_ ),
    .B(\v0/z2/z7/_012_ ),
    .Y(\v0/q1 [7]));
 sky130_fd_sc_hd__lpflow_inputiso1p_1 \v0/z2/z7/_067_  (.A(\v0/z2/q5 [4]),
    .SLEEP(\v0/z2/q4 [4]),
    .X(\v0/z2/z7/_013_ ));
 sky130_fd_sc_hd__and2_0 \v0/z2/z7/_068_  (.A(\v0/z2/q5 [4]),
    .B(\v0/z2/q4 [4]),
    .X(\v0/z2/z7/_014_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z2/z7/_069_  (.A(\v0/z2/q5 [4]),
    .B(\v0/z2/q4 [4]),
    .Y(\v0/z2/z7/_015_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z2/z7/_070_  (.A(\v0/z2/z7/_013_ ),
    .B(\v0/z2/z7/_015_ ),
    .Y(\v0/z2/z7/_016_ ));
 sky130_fd_sc_hd__o221a_1 \v0/z2/z7/_071_  (.A1(\v0/z2/q5 [3]),
    .A2(\v0/z2/q4 [3]),
    .B1(\v0/z2/z7/_003_ ),
    .B2(\v0/z2/z7/_005_ ),
    .C1(\v0/z2/z7/_004_ ),
    .X(\v0/z2/z7/_017_ ));
 sky130_fd_sc_hd__a21oi_1 \v0/z2/z7/_072_  (.A1(\v0/z2/z7/_009_ ),
    .A2(\v0/z2/z7/_012_ ),
    .B1(\v0/z2/z7/_008_ ),
    .Y(\v0/z2/z7/_018_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z2/z7/_073_  (.A(\v0/z2/z7/_016_ ),
    .B(\v0/z2/z7/_018_ ),
    .Y(\v0/q1 [8]));
 sky130_fd_sc_hd__lpflow_inputiso1p_1 \v0/z2/z7/_074_  (.A(\v0/z2/q5 [5]),
    .SLEEP(\v0/z2/q4 [5]),
    .X(\v0/z2/z7/_019_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z2/z7/_075_  (.A(\v0/z2/q5 [5]),
    .B(\v0/z2/q4 [5]),
    .Y(\v0/z2/z7/_020_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z2/z7/_076_  (.A(\v0/z2/z7/_019_ ),
    .B(\v0/z2/z7/_020_ ),
    .Y(\v0/z2/z7/_021_ ));
 sky130_fd_sc_hd__o21ai_0 \v0/z2/z7/_077_  (.A1(\v0/z2/z7/_014_ ),
    .A2(\v0/z2/z7/_018_ ),
    .B1(\v0/z2/z7/_013_ ),
    .Y(\v0/z2/z7/_022_ ));
 sky130_fd_sc_hd__xor2_1 \v0/z2/z7/_078_  (.A(\v0/z2/z7/_021_ ),
    .B(\v0/z2/z7/_022_ ),
    .X(\v0/q1 [9]));
 sky130_fd_sc_hd__nor2_1 \v0/z2/z7/_079_  (.A(\v0/z2/q5 [6]),
    .B(\v0/z2/q4 [6]),
    .Y(\v0/z2/z7/_023_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z2/z7/_080_  (.A(\v0/z2/q5 [6]),
    .B(\v0/z2/q4 [6]),
    .Y(\v0/z2/z7/_024_ ));
 sky130_fd_sc_hd__nor2b_1 \v0/z2/z7/_081_  (.A(\v0/z2/z7/_023_ ),
    .B_N(\v0/z2/z7/_024_ ),
    .Y(\v0/z2/z7/_025_ ));
 sky130_fd_sc_hd__o311ai_0 \v0/z2/z7/_082_  (.A1(\v0/z2/z7/_010_ ),
    .A2(\v0/z2/z7/_014_ ),
    .A3(\v0/z2/z7/_017_ ),
    .B1(\v0/z2/z7/_019_ ),
    .C1(\v0/z2/z7/_013_ ),
    .Y(\v0/z2/z7/_026_ ));
 sky130_fd_sc_hd__and2_0 \v0/z2/z7/_083_  (.A(\v0/z2/z7/_020_ ),
    .B(\v0/z2/z7/_026_ ),
    .X(\v0/z2/z7/_027_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z2/z7/_084_  (.A(\v0/z2/z7/_025_ ),
    .B(\v0/z2/z7/_027_ ),
    .Y(\v0/q1 [10]));
 sky130_fd_sc_hd__nor2_1 \v0/z2/z7/_085_  (.A(\v0/z2/q5 [7]),
    .B(\v0/z2/q4 [7]),
    .Y(\v0/z2/z7/_028_ ));
 sky130_fd_sc_hd__and2_0 \v0/z2/z7/_086_  (.A(\v0/z2/q5 [7]),
    .B(\v0/z2/q4 [7]),
    .X(\v0/z2/z7/_029_ ));
 sky130_fd_sc_hd__nor2_1 \v0/z2/z7/_087_  (.A(\v0/z2/z7/_028_ ),
    .B(\v0/z2/z7/_029_ ),
    .Y(\v0/z2/z7/_030_ ));
 sky130_fd_sc_hd__a21oi_1 \v0/z2/z7/_088_  (.A1(\v0/z2/z7/_024_ ),
    .A2(\v0/z2/z7/_027_ ),
    .B1(\v0/z2/z7/_023_ ),
    .Y(\v0/z2/z7/_031_ ));
 sky130_fd_sc_hd__xor2_1 \v0/z2/z7/_089_  (.A(\v0/z2/z7/_030_ ),
    .B(\v0/z2/z7/_031_ ),
    .X(\v0/q1 [11]));
 sky130_fd_sc_hd__lpflow_inputiso1p_1 \v0/z2/z7/_090_  (.A(\v0/z2/q5 [8]),
    .SLEEP(\v0/z2/_14_ ),
    .X(\v0/z2/z7/_032_ ));
 sky130_fd_sc_hd__and2_0 \v0/z2/z7/_091_  (.A(\v0/z2/q5 [8]),
    .B(\v0/z2/_14_ ),
    .X(\v0/z2/z7/_033_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z2/z7/_092_  (.A(\v0/z2/q5 [8]),
    .B(\v0/z2/_14_ ),
    .Y(\v0/z2/z7/_034_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z2/z7/_093_  (.A(\v0/z2/z7/_032_ ),
    .B(\v0/z2/z7/_034_ ),
    .Y(\v0/z2/z7/_035_ ));
 sky130_fd_sc_hd__a311oi_1 \v0/z2/z7/_094_  (.A1(\v0/z2/z7/_020_ ),
    .A2(\v0/z2/z7/_024_ ),
    .A3(\v0/z2/z7/_026_ ),
    .B1(\v0/z2/z7/_028_ ),
    .C1(\v0/z2/z7/_023_ ),
    .Y(\v0/z2/z7/_036_ ));
 sky130_fd_sc_hd__lpflow_inputiso1p_1 \v0/z2/z7/_095_  (.A(\v0/z2/z7/_029_ ),
    .SLEEP(\v0/z2/z7/_036_ ),
    .X(\v0/z2/z7/_037_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z2/z7/_096_  (.A(\v0/z2/z7/_035_ ),
    .B(\v0/z2/z7/_037_ ),
    .Y(\v0/q1 [12]));
 sky130_fd_sc_hd__lpflow_inputiso1p_1 \v0/z2/z7/_097_  (.A(\v0/z2/q5 [9]),
    .SLEEP(\v0/z2/_15_ ),
    .X(\v0/z2/z7/_038_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z2/z7/_098_  (.A(\v0/z2/q5 [9]),
    .B(\v0/z2/_15_ ),
    .Y(\v0/z2/z7/_039_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z2/z7/_099_  (.A(\v0/z2/z7/_038_ ),
    .B(\v0/z2/z7/_039_ ),
    .Y(\v0/z2/z7/_040_ ));
 sky130_fd_sc_hd__o21ai_0 \v0/z2/z7/_100_  (.A1(\v0/z2/z7/_033_ ),
    .A2(\v0/z2/z7/_037_ ),
    .B1(\v0/z2/z7/_032_ ),
    .Y(\v0/z2/z7/_041_ ));
 sky130_fd_sc_hd__xor2_1 \v0/z2/z7/_101_  (.A(\v0/z2/z7/_040_ ),
    .B(\v0/z2/z7/_041_ ),
    .X(\v0/q1 [13]));
 sky130_fd_sc_hd__nor2_1 \v0/z2/z7/_102_  (.A(\v0/z2/q5 [10]),
    .B(\v0/z2/_16_ ),
    .Y(\v0/z2/z7/_042_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z2/z7/_103_  (.A(\v0/z2/q5 [10]),
    .B(\v0/z2/_16_ ),
    .Y(\v0/z2/z7/_043_ ));
 sky130_fd_sc_hd__nand2b_1 \v0/z2/z7/_104_  (.A_N(\v0/z2/z7/_042_ ),
    .B(\v0/z2/z7/_043_ ),
    .Y(\v0/z2/z7/_044_ ));
 sky130_fd_sc_hd__o311ai_0 \v0/z2/z7/_105_  (.A1(\v0/z2/z7/_029_ ),
    .A2(\v0/z2/z7/_033_ ),
    .A3(\v0/z2/z7/_036_ ),
    .B1(\v0/z2/z7/_038_ ),
    .C1(\v0/z2/z7/_032_ ),
    .Y(\v0/z2/z7/_045_ ));
 sky130_fd_sc_hd__a21oi_1 \v0/z2/z7/_106_  (.A1(\v0/z2/z7/_039_ ),
    .A2(\v0/z2/z7/_045_ ),
    .B1(\v0/z2/z7/_044_ ),
    .Y(\v0/z2/z7/_046_ ));
 sky130_fd_sc_hd__and3_1 \v0/z2/z7/_107_  (.A(\v0/z2/z7/_039_ ),
    .B(\v0/z2/z7/_044_ ),
    .C(\v0/z2/z7/_045_ ),
    .X(\v0/z2/z7/_047_ ));
 sky130_fd_sc_hd__nor2_1 \v0/z2/z7/_108_  (.A(\v0/z2/z7/_046_ ),
    .B(\v0/z2/z7/_047_ ),
    .Y(\v0/q1 [14]));
 sky130_fd_sc_hd__xnor2_1 \v0/z2/z7/_109_  (.A(\v0/z2/q5 [11]),
    .B(\v0/z2/_17_ ),
    .Y(\v0/z2/z7/_048_ ));
 sky130_fd_sc_hd__a31oi_1 \v0/z2/z7/_110_  (.A1(\v0/z2/z7/_039_ ),
    .A2(\v0/z2/z7/_043_ ),
    .A3(\v0/z2/z7/_045_ ),
    .B1(\v0/z2/z7/_042_ ),
    .Y(\v0/z2/z7/_049_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z2/z7/_111_  (.A(\v0/z2/z7/_048_ ),
    .B(\v0/z2/z7/_049_ ),
    .Y(\v0/q1 [15]));
 sky130_fd_sc_hd__maj3_1 \v0/z2/z7/_112_  (.A(\v0/z2/q5 [11]),
    .B(\v0/z2/_17_ ),
    .C(\v0/z2/z7/_049_ ),
    .X(\v0/z2/z7/Cout ));
 sky130_fd_sc_hd__conb_1 \v0/z3/_19_  (.LO(\v0/z3/_00_ ));
 sky130_fd_sc_hd__conb_1 \v0/z3/_20_  (.LO(\v0/z3/_01_ ));
 sky130_fd_sc_hd__conb_1 \v0/z3/_21_  (.LO(\v0/z3/_02_ ));
 sky130_fd_sc_hd__conb_1 \v0/z3/_22_  (.LO(\v0/z3/_03_ ));
 sky130_fd_sc_hd__conb_1 \v0/z3/_23_  (.LO(\v0/z3/_04_ ));
 sky130_fd_sc_hd__conb_1 \v0/z3/_24_  (.LO(\v0/z3/_05_ ));
 sky130_fd_sc_hd__conb_1 \v0/z3/_25_  (.LO(\v0/z3/_06_ ));
 sky130_fd_sc_hd__conb_1 \v0/z3/_26_  (.LO(\v0/z3/_07_ ));
 sky130_fd_sc_hd__conb_1 \v0/z3/_27_  (.LO(\v0/z3/_08_ ));
 sky130_fd_sc_hd__conb_1 \v0/z3/_28_  (.LO(\v0/z3/_09_ ));
 sky130_fd_sc_hd__conb_1 \v0/z3/_29_  (.LO(\v0/z3/_10_ ));
 sky130_fd_sc_hd__conb_1 \v0/z3/_30_  (.LO(\v0/z3/_11_ ));
 sky130_fd_sc_hd__conb_1 \v0/z3/_31_  (.LO(\v0/z3/_12_ ));
 sky130_fd_sc_hd__conb_1 \v0/z3/_32_  (.LO(\v0/z3/_13_ ));
 sky130_fd_sc_hd__conb_1 \v0/z3/_33_  (.LO(\v0/z3/_14_ ));
 sky130_fd_sc_hd__conb_1 \v0/z3/_34_  (.LO(\v0/z3/_15_ ));
 sky130_fd_sc_hd__conb_1 \v0/z3/_35_  (.LO(\v0/z3/_16_ ));
 sky130_fd_sc_hd__conb_1 \v0/z3/_36_  (.LO(\v0/z3/_17_ ));
 sky130_fd_sc_hd__conb_1 \v0/z3/_37_  (.LO(\v0/z3/_18_ ));
 sky130_fd_sc_hd__conb_1 \v0/z3/z1/_11_  (.LO(\v0/z3/z1/_00_ ));
 sky130_fd_sc_hd__conb_1 \v0/z3/z1/_12_  (.LO(\v0/z3/z1/_01_ ));
 sky130_fd_sc_hd__conb_1 \v0/z3/z1/_13_  (.LO(\v0/z3/z1/_02_ ));
 sky130_fd_sc_hd__conb_1 \v0/z3/z1/_14_  (.LO(\v0/z3/z1/_03_ ));
 sky130_fd_sc_hd__conb_1 \v0/z3/z1/_15_  (.LO(\v0/z3/z1/_04_ ));
 sky130_fd_sc_hd__conb_1 \v0/z3/z1/_16_  (.LO(\v0/z3/z1/_05_ ));
 sky130_fd_sc_hd__conb_1 \v0/z3/z1/_17_  (.LO(\v0/z3/z1/_06_ ));
 sky130_fd_sc_hd__conb_1 \v0/z3/z1/_18_  (.LO(\v0/z3/z1/_07_ ));
 sky130_fd_sc_hd__conb_1 \v0/z3/z1/_19_  (.LO(\v0/z3/z1/_08_ ));
 sky130_fd_sc_hd__conb_1 \v0/z3/z1/_20_  (.LO(\v0/z3/z1/_09_ ));
 sky130_fd_sc_hd__conb_1 \v0/z3/z1/_21_  (.LO(\v0/z3/z1/_10_ ));
 sky130_fd_sc_hd__and2_0 \v0/z3/z1/z1/_0_  (.A(abs_b[8]),
    .B(a[0]),
    .X(\v0/q2 [0]));
 sky130_fd_sc_hd__and2_0 \v0/z3/z1/z1/_1_  (.A(abs_b[8]),
    .B(abs_a[1]),
    .X(\v0/z3/z1/z1/temp [0]));
 sky130_fd_sc_hd__and2_0 \v0/z3/z1/z1/_2_  (.A(a[0]),
    .B(abs_b[9]),
    .X(\v0/z3/z1/z1/temp [1]));
 sky130_fd_sc_hd__and2_0 \v0/z3/z1/z1/_3_  (.A(abs_a[1]),
    .B(abs_b[9]),
    .X(\v0/z3/z1/z1/temp [2]));
 sky130_fd_sc_hd__and2_0 \v0/z3/z1/z1/z1/_0_  (.A(\v0/z3/z1/z1/temp [1]),
    .B(\v0/z3/z1/z1/temp [0]),
    .X(\v0/z3/z1/z1/temp [3]));
 sky130_fd_sc_hd__xor2_1 \v0/z3/z1/z1/z1/_1_  (.A(\v0/z3/z1/z1/temp [1]),
    .B(\v0/z3/z1/z1/temp [0]),
    .X(\v0/q2 [1]));
 sky130_fd_sc_hd__and2_0 \v0/z3/z1/z1/z2/_0_  (.A(\v0/z3/z1/z1/temp [3]),
    .B(\v0/z3/z1/z1/temp [2]),
    .X(\v0/z3/z1/q0 [3]));
 sky130_fd_sc_hd__xor2_1 \v0/z3/z1/z1/z2/_1_  (.A(\v0/z3/z1/z1/temp [3]),
    .B(\v0/z3/z1/z1/temp [2]),
    .X(\v0/z3/z1/q0 [2]));
 sky130_fd_sc_hd__and2_0 \v0/z3/z1/z2/_0_  (.A(abs_b[8]),
    .B(abs_a[2]),
    .X(\v0/z3/z1/q1 [0]));
 sky130_fd_sc_hd__and2_0 \v0/z3/z1/z2/_1_  (.A(abs_b[8]),
    .B(abs_a[3]),
    .X(\v0/z3/z1/z2/temp [0]));
 sky130_fd_sc_hd__and2_0 \v0/z3/z1/z2/_2_  (.A(abs_a[2]),
    .B(abs_b[9]),
    .X(\v0/z3/z1/z2/temp [1]));
 sky130_fd_sc_hd__and2_0 \v0/z3/z1/z2/_3_  (.A(abs_a[3]),
    .B(abs_b[9]),
    .X(\v0/z3/z1/z2/temp [2]));
 sky130_fd_sc_hd__and2_0 \v0/z3/z1/z2/z1/_0_  (.A(\v0/z3/z1/z2/temp [1]),
    .B(\v0/z3/z1/z2/temp [0]),
    .X(\v0/z3/z1/z2/temp [3]));
 sky130_fd_sc_hd__xor2_1 \v0/z3/z1/z2/z1/_1_  (.A(\v0/z3/z1/z2/temp [1]),
    .B(\v0/z3/z1/z2/temp [0]),
    .X(\v0/z3/z1/q1 [1]));
 sky130_fd_sc_hd__and2_0 \v0/z3/z1/z2/z2/_0_  (.A(\v0/z3/z1/z2/temp [3]),
    .B(\v0/z3/z1/z2/temp [2]),
    .X(\v0/z3/z1/q1 [3]));
 sky130_fd_sc_hd__xor2_1 \v0/z3/z1/z2/z2/_1_  (.A(\v0/z3/z1/z2/temp [3]),
    .B(\v0/z3/z1/z2/temp [2]),
    .X(\v0/z3/z1/q1 [2]));
 sky130_fd_sc_hd__and2_0 \v0/z3/z1/z3/_0_  (.A(abs_b[10]),
    .B(a[0]),
    .X(\v0/z3/z1/q2 [0]));
 sky130_fd_sc_hd__and2_0 \v0/z3/z1/z3/_1_  (.A(abs_b[10]),
    .B(abs_a[1]),
    .X(\v0/z3/z1/z3/temp [0]));
 sky130_fd_sc_hd__and2_0 \v0/z3/z1/z3/_2_  (.A(a[0]),
    .B(abs_b[11]),
    .X(\v0/z3/z1/z3/temp [1]));
 sky130_fd_sc_hd__and2_0 \v0/z3/z1/z3/_3_  (.A(abs_a[1]),
    .B(abs_b[11]),
    .X(\v0/z3/z1/z3/temp [2]));
 sky130_fd_sc_hd__and2_0 \v0/z3/z1/z3/z1/_0_  (.A(\v0/z3/z1/z3/temp [1]),
    .B(\v0/z3/z1/z3/temp [0]),
    .X(\v0/z3/z1/z3/temp [3]));
 sky130_fd_sc_hd__xor2_1 \v0/z3/z1/z3/z1/_1_  (.A(\v0/z3/z1/z3/temp [1]),
    .B(\v0/z3/z1/z3/temp [0]),
    .X(\v0/z3/z1/q2 [1]));
 sky130_fd_sc_hd__and2_0 \v0/z3/z1/z3/z2/_0_  (.A(\v0/z3/z1/z3/temp [3]),
    .B(\v0/z3/z1/z3/temp [2]),
    .X(\v0/z3/z1/q2 [3]));
 sky130_fd_sc_hd__xor2_1 \v0/z3/z1/z3/z2/_1_  (.A(\v0/z3/z1/z3/temp [3]),
    .B(\v0/z3/z1/z3/temp [2]),
    .X(\v0/z3/z1/q2 [2]));
 sky130_fd_sc_hd__and2_0 \v0/z3/z1/z4/_0_  (.A(abs_b[10]),
    .B(abs_a[2]),
    .X(\v0/z3/z1/q3 [0]));
 sky130_fd_sc_hd__and2_0 \v0/z3/z1/z4/_1_  (.A(abs_b[10]),
    .B(abs_a[3]),
    .X(\v0/z3/z1/z4/temp [0]));
 sky130_fd_sc_hd__and2_0 \v0/z3/z1/z4/_2_  (.A(abs_a[2]),
    .B(abs_b[11]),
    .X(\v0/z3/z1/z4/temp [1]));
 sky130_fd_sc_hd__and2_0 \v0/z3/z1/z4/_3_  (.A(abs_a[3]),
    .B(abs_b[11]),
    .X(\v0/z3/z1/z4/temp [2]));
 sky130_fd_sc_hd__and2_0 \v0/z3/z1/z4/z1/_0_  (.A(\v0/z3/z1/z4/temp [1]),
    .B(\v0/z3/z1/z4/temp [0]),
    .X(\v0/z3/z1/z4/temp [3]));
 sky130_fd_sc_hd__xor2_1 \v0/z3/z1/z4/z1/_1_  (.A(\v0/z3/z1/z4/temp [1]),
    .B(\v0/z3/z1/z4/temp [0]),
    .X(\v0/z3/z1/q3 [1]));
 sky130_fd_sc_hd__and2_0 \v0/z3/z1/z4/z2/_0_  (.A(\v0/z3/z1/z4/temp [3]),
    .B(\v0/z3/z1/z4/temp [2]),
    .X(\v0/z3/z1/q3 [3]));
 sky130_fd_sc_hd__xor2_1 \v0/z3/z1/z4/z2/_1_  (.A(\v0/z3/z1/z4/temp [3]),
    .B(\v0/z3/z1/z4/temp [2]),
    .X(\v0/z3/z1/q3 [2]));
 sky130_fd_sc_hd__xnor2_1 \v0/z3/z1/z5/_07_  (.A(\v0/z3/z1/q0 [2]),
    .B(\v0/z3/z1/q1 [0]),
    .Y(\v0/z3/z1/z5/_00_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z3/z1/z5/_08_  (.A(\v0/z3/z1/_02_ ),
    .B(\v0/z3/z1/z5/_00_ ),
    .Y(\v0/z3/z1/q4 [0]));
 sky130_fd_sc_hd__maj3_1 \v0/z3/z1/z5/_09_  (.A(\v0/z3/z1/q0 [2]),
    .B(\v0/z3/z1/q1 [0]),
    .C(\v0/z3/z1/_02_ ),
    .X(\v0/z3/z1/z5/_01_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z3/z1/z5/_10_  (.A(\v0/z3/z1/q0 [3]),
    .B(\v0/z3/z1/q1 [1]),
    .Y(\v0/z3/z1/z5/_02_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z3/z1/z5/_11_  (.A(\v0/z3/z1/z5/_01_ ),
    .B(\v0/z3/z1/z5/_02_ ),
    .Y(\v0/z3/z1/q4 [1]));
 sky130_fd_sc_hd__maj3_1 \v0/z3/z1/z5/_12_  (.A(\v0/z3/z1/q0 [3]),
    .B(\v0/z3/z1/q1 [1]),
    .C(\v0/z3/z1/z5/_01_ ),
    .X(\v0/z3/z1/z5/_03_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z3/z1/z5/_13_  (.A(\v0/z3/z1/_00_ ),
    .B(\v0/z3/z1/q1 [2]),
    .Y(\v0/z3/z1/z5/_04_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z3/z1/z5/_14_  (.A(\v0/z3/z1/z5/_03_ ),
    .B(\v0/z3/z1/z5/_04_ ),
    .Y(\v0/z3/z1/q4 [2]));
 sky130_fd_sc_hd__maj3_1 \v0/z3/z1/z5/_15_  (.A(\v0/z3/z1/_00_ ),
    .B(\v0/z3/z1/q1 [2]),
    .C(\v0/z3/z1/z5/_03_ ),
    .X(\v0/z3/z1/z5/_05_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z3/z1/z5/_16_  (.A(\v0/z3/z1/_01_ ),
    .B(\v0/z3/z1/q1 [3]),
    .Y(\v0/z3/z1/z5/_06_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z3/z1/z5/_17_  (.A(\v0/z3/z1/z5/_05_ ),
    .B(\v0/z3/z1/z5/_06_ ),
    .Y(\v0/z3/z1/q4 [3]));
 sky130_fd_sc_hd__maj3_1 \v0/z3/z1/z5/_18_  (.A(\v0/z3/z1/_01_ ),
    .B(\v0/z3/z1/q1 [3]),
    .C(\v0/z3/z1/z5/_05_ ),
    .X(\v0/z3/z1/z5/Cout ));
 sky130_fd_sc_hd__xnor2_1 \v0/z3/z1/z6/_19_  (.A(\v0/z3/z1/_05_ ),
    .B(\v0/z3/z1/q2 [0]),
    .Y(\v0/z3/z1/z6/_00_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z3/z1/z6/_20_  (.A(\v0/z3/z1/_07_ ),
    .B(\v0/z3/z1/z6/_00_ ),
    .Y(\v0/z3/z1/q5 [0]));
 sky130_fd_sc_hd__maj3_1 \v0/z3/z1/z6/_21_  (.A(\v0/z3/z1/_05_ ),
    .B(\v0/z3/z1/q2 [0]),
    .C(\v0/z3/z1/_07_ ),
    .X(\v0/z3/z1/z6/_01_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z3/z1/z6/_22_  (.A(\v0/z3/z1/_06_ ),
    .B(\v0/z3/z1/q2 [1]),
    .Y(\v0/z3/z1/z6/_02_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z3/z1/z6/_23_  (.A(\v0/z3/z1/z6/_01_ ),
    .B(\v0/z3/z1/z6/_02_ ),
    .Y(\v0/z3/z1/q5 [1]));
 sky130_fd_sc_hd__maj3_1 \v0/z3/z1/z6/_24_  (.A(\v0/z3/z1/_06_ ),
    .B(\v0/z3/z1/q2 [1]),
    .C(\v0/z3/z1/z6/_01_ ),
    .X(\v0/z3/z1/z6/_03_ ));
 sky130_fd_sc_hd__lpflow_inputiso1p_1 \v0/z3/z1/z6/_25_  (.A(\v0/z3/z1/q3 [0]),
    .SLEEP(\v0/z3/z1/q2 [2]),
    .X(\v0/z3/z1/z6/_04_ ));
 sky130_fd_sc_hd__and2_0 \v0/z3/z1/z6/_26_  (.A(\v0/z3/z1/q3 [0]),
    .B(\v0/z3/z1/q2 [2]),
    .X(\v0/z3/z1/z6/_05_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z3/z1/z6/_27_  (.A(\v0/z3/z1/q3 [0]),
    .B(\v0/z3/z1/q2 [2]),
    .Y(\v0/z3/z1/z6/_06_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z3/z1/z6/_28_  (.A(\v0/z3/z1/z6/_04_ ),
    .B(\v0/z3/z1/z6/_06_ ),
    .Y(\v0/z3/z1/z6/_07_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z3/z1/z6/_29_  (.A(\v0/z3/z1/z6/_03_ ),
    .B(\v0/z3/z1/z6/_07_ ),
    .Y(\v0/z3/z1/q5 [2]));
 sky130_fd_sc_hd__nand2_1 \v0/z3/z1/z6/_30_  (.A(\v0/z3/z1/q3 [1]),
    .B(\v0/z3/z1/q2 [3]),
    .Y(\v0/z3/z1/z6/_08_ ));
 sky130_fd_sc_hd__xor2_1 \v0/z3/z1/z6/_31_  (.A(\v0/z3/z1/q3 [1]),
    .B(\v0/z3/z1/q2 [3]),
    .X(\v0/z3/z1/z6/_09_ ));
 sky130_fd_sc_hd__o21ai_0 \v0/z3/z1/z6/_32_  (.A1(\v0/z3/z1/z6/_03_ ),
    .A2(\v0/z3/z1/z6/_05_ ),
    .B1(\v0/z3/z1/z6/_04_ ),
    .Y(\v0/z3/z1/z6/_10_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z3/z1/z6/_33_  (.A(\v0/z3/z1/z6/_09_ ),
    .B(\v0/z3/z1/z6/_10_ ),
    .Y(\v0/z3/z1/q5 [3]));
 sky130_fd_sc_hd__nor2_1 \v0/z3/z1/z6/_34_  (.A(\v0/z3/z1/q3 [2]),
    .B(\v0/z3/z1/_03_ ),
    .Y(\v0/z3/z1/z6/_11_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z3/z1/z6/_35_  (.A(\v0/z3/z1/q3 [2]),
    .B(\v0/z3/z1/_03_ ),
    .Y(\v0/z3/z1/z6/_12_ ));
 sky130_fd_sc_hd__nand2b_1 \v0/z3/z1/z6/_36_  (.A_N(\v0/z3/z1/z6/_11_ ),
    .B(\v0/z3/z1/z6/_12_ ),
    .Y(\v0/z3/z1/z6/_13_ ));
 sky130_fd_sc_hd__o221ai_1 \v0/z3/z1/z6/_37_  (.A1(\v0/z3/z1/q3 [1]),
    .A2(\v0/z3/z1/q2 [3]),
    .B1(\v0/z3/z1/z6/_03_ ),
    .B2(\v0/z3/z1/z6/_05_ ),
    .C1(\v0/z3/z1/z6/_04_ ),
    .Y(\v0/z3/z1/z6/_14_ ));
 sky130_fd_sc_hd__a21oi_1 \v0/z3/z1/z6/_38_  (.A1(\v0/z3/z1/z6/_08_ ),
    .A2(\v0/z3/z1/z6/_14_ ),
    .B1(\v0/z3/z1/z6/_13_ ),
    .Y(\v0/z3/z1/z6/_15_ ));
 sky130_fd_sc_hd__and3_1 \v0/z3/z1/z6/_39_  (.A(\v0/z3/z1/z6/_08_ ),
    .B(\v0/z3/z1/z6/_13_ ),
    .C(\v0/z3/z1/z6/_14_ ),
    .X(\v0/z3/z1/z6/_16_ ));
 sky130_fd_sc_hd__nor2_1 \v0/z3/z1/z6/_40_  (.A(\v0/z3/z1/z6/_15_ ),
    .B(\v0/z3/z1/z6/_16_ ),
    .Y(\v0/z3/z1/q5 [4]));
 sky130_fd_sc_hd__xnor2_1 \v0/z3/z1/z6/_41_  (.A(\v0/z3/z1/q3 [3]),
    .B(\v0/z3/z1/_04_ ),
    .Y(\v0/z3/z1/z6/_17_ ));
 sky130_fd_sc_hd__a31oi_1 \v0/z3/z1/z6/_42_  (.A1(\v0/z3/z1/z6/_08_ ),
    .A2(\v0/z3/z1/z6/_12_ ),
    .A3(\v0/z3/z1/z6/_14_ ),
    .B1(\v0/z3/z1/z6/_11_ ),
    .Y(\v0/z3/z1/z6/_18_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z3/z1/z6/_43_  (.A(\v0/z3/z1/z6/_17_ ),
    .B(\v0/z3/z1/z6/_18_ ),
    .Y(\v0/z3/z1/q5 [5]));
 sky130_fd_sc_hd__maj3_1 \v0/z3/z1/z6/_44_  (.A(\v0/z3/z1/q3 [3]),
    .B(\v0/z3/z1/_04_ ),
    .C(\v0/z3/z1/z6/_18_ ),
    .X(\v0/z3/z1/z6/Cout ));
 sky130_fd_sc_hd__xnor2_1 \v0/z3/z1/z7/_19_  (.A(\v0/z3/z1/q5 [0]),
    .B(\v0/z3/z1/q4 [0]),
    .Y(\v0/z3/z1/z7/_00_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z3/z1/z7/_20_  (.A(\v0/z3/z1/_10_ ),
    .B(\v0/z3/z1/z7/_00_ ),
    .Y(\v0/q2 [2]));
 sky130_fd_sc_hd__maj3_1 \v0/z3/z1/z7/_21_  (.A(\v0/z3/z1/q5 [0]),
    .B(\v0/z3/z1/q4 [0]),
    .C(\v0/z3/z1/_10_ ),
    .X(\v0/z3/z1/z7/_01_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z3/z1/z7/_22_  (.A(\v0/z3/z1/q5 [1]),
    .B(\v0/z3/z1/q4 [1]),
    .Y(\v0/z3/z1/z7/_02_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z3/z1/z7/_23_  (.A(\v0/z3/z1/z7/_01_ ),
    .B(\v0/z3/z1/z7/_02_ ),
    .Y(\v0/q2 [3]));
 sky130_fd_sc_hd__maj3_1 \v0/z3/z1/z7/_24_  (.A(\v0/z3/z1/q5 [1]),
    .B(\v0/z3/z1/q4 [1]),
    .C(\v0/z3/z1/z7/_01_ ),
    .X(\v0/z3/z1/z7/_03_ ));
 sky130_fd_sc_hd__lpflow_inputiso1p_1 \v0/z3/z1/z7/_25_  (.A(\v0/z3/z1/q5 [2]),
    .SLEEP(\v0/z3/z1/q4 [2]),
    .X(\v0/z3/z1/z7/_04_ ));
 sky130_fd_sc_hd__and2_0 \v0/z3/z1/z7/_26_  (.A(\v0/z3/z1/q5 [2]),
    .B(\v0/z3/z1/q4 [2]),
    .X(\v0/z3/z1/z7/_05_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z3/z1/z7/_27_  (.A(\v0/z3/z1/q5 [2]),
    .B(\v0/z3/z1/q4 [2]),
    .Y(\v0/z3/z1/z7/_06_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z3/z1/z7/_28_  (.A(\v0/z3/z1/z7/_04_ ),
    .B(\v0/z3/z1/z7/_06_ ),
    .Y(\v0/z3/z1/z7/_07_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z3/z1/z7/_29_  (.A(\v0/z3/z1/z7/_03_ ),
    .B(\v0/z3/z1/z7/_07_ ),
    .Y(\v0/z3/q0 [4]));
 sky130_fd_sc_hd__nand2_1 \v0/z3/z1/z7/_30_  (.A(\v0/z3/z1/q5 [3]),
    .B(\v0/z3/z1/q4 [3]),
    .Y(\v0/z3/z1/z7/_08_ ));
 sky130_fd_sc_hd__xor2_1 \v0/z3/z1/z7/_31_  (.A(\v0/z3/z1/q5 [3]),
    .B(\v0/z3/z1/q4 [3]),
    .X(\v0/z3/z1/z7/_09_ ));
 sky130_fd_sc_hd__o21ai_0 \v0/z3/z1/z7/_32_  (.A1(\v0/z3/z1/z7/_03_ ),
    .A2(\v0/z3/z1/z7/_05_ ),
    .B1(\v0/z3/z1/z7/_04_ ),
    .Y(\v0/z3/z1/z7/_10_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z3/z1/z7/_33_  (.A(\v0/z3/z1/z7/_09_ ),
    .B(\v0/z3/z1/z7/_10_ ),
    .Y(\v0/z3/q0 [5]));
 sky130_fd_sc_hd__nor2_1 \v0/z3/z1/z7/_34_  (.A(\v0/z3/z1/q5 [4]),
    .B(\v0/z3/z1/_08_ ),
    .Y(\v0/z3/z1/z7/_11_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z3/z1/z7/_35_  (.A(\v0/z3/z1/q5 [4]),
    .B(\v0/z3/z1/_08_ ),
    .Y(\v0/z3/z1/z7/_12_ ));
 sky130_fd_sc_hd__nand2b_1 \v0/z3/z1/z7/_36_  (.A_N(\v0/z3/z1/z7/_11_ ),
    .B(\v0/z3/z1/z7/_12_ ),
    .Y(\v0/z3/z1/z7/_13_ ));
 sky130_fd_sc_hd__o221ai_1 \v0/z3/z1/z7/_37_  (.A1(\v0/z3/z1/q5 [3]),
    .A2(\v0/z3/z1/q4 [3]),
    .B1(\v0/z3/z1/z7/_03_ ),
    .B2(\v0/z3/z1/z7/_05_ ),
    .C1(\v0/z3/z1/z7/_04_ ),
    .Y(\v0/z3/z1/z7/_14_ ));
 sky130_fd_sc_hd__a21oi_1 \v0/z3/z1/z7/_38_  (.A1(\v0/z3/z1/z7/_08_ ),
    .A2(\v0/z3/z1/z7/_14_ ),
    .B1(\v0/z3/z1/z7/_13_ ),
    .Y(\v0/z3/z1/z7/_15_ ));
 sky130_fd_sc_hd__and3_1 \v0/z3/z1/z7/_39_  (.A(\v0/z3/z1/z7/_08_ ),
    .B(\v0/z3/z1/z7/_13_ ),
    .C(\v0/z3/z1/z7/_14_ ),
    .X(\v0/z3/z1/z7/_16_ ));
 sky130_fd_sc_hd__nor2_1 \v0/z3/z1/z7/_40_  (.A(\v0/z3/z1/z7/_15_ ),
    .B(\v0/z3/z1/z7/_16_ ),
    .Y(\v0/z3/q0 [6]));
 sky130_fd_sc_hd__xnor2_1 \v0/z3/z1/z7/_41_  (.A(\v0/z3/z1/q5 [5]),
    .B(\v0/z3/z1/_09_ ),
    .Y(\v0/z3/z1/z7/_17_ ));
 sky130_fd_sc_hd__a31oi_1 \v0/z3/z1/z7/_42_  (.A1(\v0/z3/z1/z7/_08_ ),
    .A2(\v0/z3/z1/z7/_12_ ),
    .A3(\v0/z3/z1/z7/_14_ ),
    .B1(\v0/z3/z1/z7/_11_ ),
    .Y(\v0/z3/z1/z7/_18_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z3/z1/z7/_43_  (.A(\v0/z3/z1/z7/_17_ ),
    .B(\v0/z3/z1/z7/_18_ ),
    .Y(\v0/z3/q0 [7]));
 sky130_fd_sc_hd__maj3_1 \v0/z3/z1/z7/_44_  (.A(\v0/z3/z1/q5 [5]),
    .B(\v0/z3/z1/_09_ ),
    .C(\v0/z3/z1/z7/_18_ ),
    .X(\v0/z3/z1/z7/Cout ));
 sky130_fd_sc_hd__conb_1 \v0/z3/z2/_11_  (.LO(\v0/z3/z2/_00_ ));
 sky130_fd_sc_hd__conb_1 \v0/z3/z2/_12_  (.LO(\v0/z3/z2/_01_ ));
 sky130_fd_sc_hd__conb_1 \v0/z3/z2/_13_  (.LO(\v0/z3/z2/_02_ ));
 sky130_fd_sc_hd__conb_1 \v0/z3/z2/_14_  (.LO(\v0/z3/z2/_03_ ));
 sky130_fd_sc_hd__conb_1 \v0/z3/z2/_15_  (.LO(\v0/z3/z2/_04_ ));
 sky130_fd_sc_hd__conb_1 \v0/z3/z2/_16_  (.LO(\v0/z3/z2/_05_ ));
 sky130_fd_sc_hd__conb_1 \v0/z3/z2/_17_  (.LO(\v0/z3/z2/_06_ ));
 sky130_fd_sc_hd__conb_1 \v0/z3/z2/_18_  (.LO(\v0/z3/z2/_07_ ));
 sky130_fd_sc_hd__conb_1 \v0/z3/z2/_19_  (.LO(\v0/z3/z2/_08_ ));
 sky130_fd_sc_hd__conb_1 \v0/z3/z2/_20_  (.LO(\v0/z3/z2/_09_ ));
 sky130_fd_sc_hd__conb_1 \v0/z3/z2/_21_  (.LO(\v0/z3/z2/_10_ ));
 sky130_fd_sc_hd__and2_0 \v0/z3/z2/z1/_0_  (.A(abs_b[8]),
    .B(abs_a[4]),
    .X(\v0/z3/q1 [0]));
 sky130_fd_sc_hd__and2_0 \v0/z3/z2/z1/_1_  (.A(abs_b[8]),
    .B(abs_a[5]),
    .X(\v0/z3/z2/z1/temp [0]));
 sky130_fd_sc_hd__and2_0 \v0/z3/z2/z1/_2_  (.A(abs_a[4]),
    .B(abs_b[9]),
    .X(\v0/z3/z2/z1/temp [1]));
 sky130_fd_sc_hd__and2_0 \v0/z3/z2/z1/_3_  (.A(abs_a[5]),
    .B(abs_b[9]),
    .X(\v0/z3/z2/z1/temp [2]));
 sky130_fd_sc_hd__and2_0 \v0/z3/z2/z1/z1/_0_  (.A(\v0/z3/z2/z1/temp [1]),
    .B(\v0/z3/z2/z1/temp [0]),
    .X(\v0/z3/z2/z1/temp [3]));
 sky130_fd_sc_hd__xor2_1 \v0/z3/z2/z1/z1/_1_  (.A(\v0/z3/z2/z1/temp [1]),
    .B(\v0/z3/z2/z1/temp [0]),
    .X(\v0/z3/q1 [1]));
 sky130_fd_sc_hd__and2_0 \v0/z3/z2/z1/z2/_0_  (.A(\v0/z3/z2/z1/temp [3]),
    .B(\v0/z3/z2/z1/temp [2]),
    .X(\v0/z3/z2/q0 [3]));
 sky130_fd_sc_hd__xor2_1 \v0/z3/z2/z1/z2/_1_  (.A(\v0/z3/z2/z1/temp [3]),
    .B(\v0/z3/z2/z1/temp [2]),
    .X(\v0/z3/z2/q0 [2]));
 sky130_fd_sc_hd__and2_0 \v0/z3/z2/z2/_0_  (.A(abs_b[8]),
    .B(abs_a[6]),
    .X(\v0/z3/z2/q1 [0]));
 sky130_fd_sc_hd__and2_0 \v0/z3/z2/z2/_1_  (.A(abs_b[8]),
    .B(abs_a[7]),
    .X(\v0/z3/z2/z2/temp [0]));
 sky130_fd_sc_hd__and2_0 \v0/z3/z2/z2/_2_  (.A(abs_a[6]),
    .B(abs_b[9]),
    .X(\v0/z3/z2/z2/temp [1]));
 sky130_fd_sc_hd__and2_0 \v0/z3/z2/z2/_3_  (.A(abs_a[7]),
    .B(abs_b[9]),
    .X(\v0/z3/z2/z2/temp [2]));
 sky130_fd_sc_hd__and2_0 \v0/z3/z2/z2/z1/_0_  (.A(\v0/z3/z2/z2/temp [1]),
    .B(\v0/z3/z2/z2/temp [0]),
    .X(\v0/z3/z2/z2/temp [3]));
 sky130_fd_sc_hd__xor2_1 \v0/z3/z2/z2/z1/_1_  (.A(\v0/z3/z2/z2/temp [1]),
    .B(\v0/z3/z2/z2/temp [0]),
    .X(\v0/z3/z2/q1 [1]));
 sky130_fd_sc_hd__and2_0 \v0/z3/z2/z2/z2/_0_  (.A(\v0/z3/z2/z2/temp [3]),
    .B(\v0/z3/z2/z2/temp [2]),
    .X(\v0/z3/z2/q1 [3]));
 sky130_fd_sc_hd__xor2_1 \v0/z3/z2/z2/z2/_1_  (.A(\v0/z3/z2/z2/temp [3]),
    .B(\v0/z3/z2/z2/temp [2]),
    .X(\v0/z3/z2/q1 [2]));
 sky130_fd_sc_hd__and2_0 \v0/z3/z2/z3/_0_  (.A(abs_b[10]),
    .B(abs_a[4]),
    .X(\v0/z3/z2/q2 [0]));
 sky130_fd_sc_hd__and2_0 \v0/z3/z2/z3/_1_  (.A(abs_b[10]),
    .B(abs_a[5]),
    .X(\v0/z3/z2/z3/temp [0]));
 sky130_fd_sc_hd__and2_0 \v0/z3/z2/z3/_2_  (.A(abs_a[4]),
    .B(abs_b[11]),
    .X(\v0/z3/z2/z3/temp [1]));
 sky130_fd_sc_hd__and2_0 \v0/z3/z2/z3/_3_  (.A(abs_a[5]),
    .B(abs_b[11]),
    .X(\v0/z3/z2/z3/temp [2]));
 sky130_fd_sc_hd__and2_0 \v0/z3/z2/z3/z1/_0_  (.A(\v0/z3/z2/z3/temp [1]),
    .B(\v0/z3/z2/z3/temp [0]),
    .X(\v0/z3/z2/z3/temp [3]));
 sky130_fd_sc_hd__xor2_1 \v0/z3/z2/z3/z1/_1_  (.A(\v0/z3/z2/z3/temp [1]),
    .B(\v0/z3/z2/z3/temp [0]),
    .X(\v0/z3/z2/q2 [1]));
 sky130_fd_sc_hd__and2_0 \v0/z3/z2/z3/z2/_0_  (.A(\v0/z3/z2/z3/temp [3]),
    .B(\v0/z3/z2/z3/temp [2]),
    .X(\v0/z3/z2/q2 [3]));
 sky130_fd_sc_hd__xor2_1 \v0/z3/z2/z3/z2/_1_  (.A(\v0/z3/z2/z3/temp [3]),
    .B(\v0/z3/z2/z3/temp [2]),
    .X(\v0/z3/z2/q2 [2]));
 sky130_fd_sc_hd__and2_0 \v0/z3/z2/z4/_0_  (.A(abs_b[10]),
    .B(abs_a[6]),
    .X(\v0/z3/z2/q3 [0]));
 sky130_fd_sc_hd__and2_0 \v0/z3/z2/z4/_1_  (.A(abs_b[10]),
    .B(abs_a[7]),
    .X(\v0/z3/z2/z4/temp [0]));
 sky130_fd_sc_hd__and2_0 \v0/z3/z2/z4/_2_  (.A(abs_a[6]),
    .B(abs_b[11]),
    .X(\v0/z3/z2/z4/temp [1]));
 sky130_fd_sc_hd__and2_0 \v0/z3/z2/z4/_3_  (.A(abs_a[7]),
    .B(abs_b[11]),
    .X(\v0/z3/z2/z4/temp [2]));
 sky130_fd_sc_hd__and2_0 \v0/z3/z2/z4/z1/_0_  (.A(\v0/z3/z2/z4/temp [1]),
    .B(\v0/z3/z2/z4/temp [0]),
    .X(\v0/z3/z2/z4/temp [3]));
 sky130_fd_sc_hd__xor2_1 \v0/z3/z2/z4/z1/_1_  (.A(\v0/z3/z2/z4/temp [1]),
    .B(\v0/z3/z2/z4/temp [0]),
    .X(\v0/z3/z2/q3 [1]));
 sky130_fd_sc_hd__and2_0 \v0/z3/z2/z4/z2/_0_  (.A(\v0/z3/z2/z4/temp [3]),
    .B(\v0/z3/z2/z4/temp [2]),
    .X(\v0/z3/z2/q3 [3]));
 sky130_fd_sc_hd__xor2_1 \v0/z3/z2/z4/z2/_1_  (.A(\v0/z3/z2/z4/temp [3]),
    .B(\v0/z3/z2/z4/temp [2]),
    .X(\v0/z3/z2/q3 [2]));
 sky130_fd_sc_hd__xnor2_1 \v0/z3/z2/z5/_07_  (.A(\v0/z3/z2/q0 [2]),
    .B(\v0/z3/z2/q1 [0]),
    .Y(\v0/z3/z2/z5/_00_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z3/z2/z5/_08_  (.A(\v0/z3/z2/_02_ ),
    .B(\v0/z3/z2/z5/_00_ ),
    .Y(\v0/z3/z2/q4 [0]));
 sky130_fd_sc_hd__maj3_1 \v0/z3/z2/z5/_09_  (.A(\v0/z3/z2/q0 [2]),
    .B(\v0/z3/z2/q1 [0]),
    .C(\v0/z3/z2/_02_ ),
    .X(\v0/z3/z2/z5/_01_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z3/z2/z5/_10_  (.A(\v0/z3/z2/q0 [3]),
    .B(\v0/z3/z2/q1 [1]),
    .Y(\v0/z3/z2/z5/_02_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z3/z2/z5/_11_  (.A(\v0/z3/z2/z5/_01_ ),
    .B(\v0/z3/z2/z5/_02_ ),
    .Y(\v0/z3/z2/q4 [1]));
 sky130_fd_sc_hd__maj3_1 \v0/z3/z2/z5/_12_  (.A(\v0/z3/z2/q0 [3]),
    .B(\v0/z3/z2/q1 [1]),
    .C(\v0/z3/z2/z5/_01_ ),
    .X(\v0/z3/z2/z5/_03_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z3/z2/z5/_13_  (.A(\v0/z3/z2/_00_ ),
    .B(\v0/z3/z2/q1 [2]),
    .Y(\v0/z3/z2/z5/_04_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z3/z2/z5/_14_  (.A(\v0/z3/z2/z5/_03_ ),
    .B(\v0/z3/z2/z5/_04_ ),
    .Y(\v0/z3/z2/q4 [2]));
 sky130_fd_sc_hd__maj3_1 \v0/z3/z2/z5/_15_  (.A(\v0/z3/z2/_00_ ),
    .B(\v0/z3/z2/q1 [2]),
    .C(\v0/z3/z2/z5/_03_ ),
    .X(\v0/z3/z2/z5/_05_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z3/z2/z5/_16_  (.A(\v0/z3/z2/_01_ ),
    .B(\v0/z3/z2/q1 [3]),
    .Y(\v0/z3/z2/z5/_06_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z3/z2/z5/_17_  (.A(\v0/z3/z2/z5/_05_ ),
    .B(\v0/z3/z2/z5/_06_ ),
    .Y(\v0/z3/z2/q4 [3]));
 sky130_fd_sc_hd__maj3_1 \v0/z3/z2/z5/_18_  (.A(\v0/z3/z2/_01_ ),
    .B(\v0/z3/z2/q1 [3]),
    .C(\v0/z3/z2/z5/_05_ ),
    .X(\v0/z3/z2/z5/Cout ));
 sky130_fd_sc_hd__xnor2_1 \v0/z3/z2/z6/_19_  (.A(\v0/z3/z2/_05_ ),
    .B(\v0/z3/z2/q2 [0]),
    .Y(\v0/z3/z2/z6/_00_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z3/z2/z6/_20_  (.A(\v0/z3/z2/_07_ ),
    .B(\v0/z3/z2/z6/_00_ ),
    .Y(\v0/z3/z2/q5 [0]));
 sky130_fd_sc_hd__maj3_1 \v0/z3/z2/z6/_21_  (.A(\v0/z3/z2/_05_ ),
    .B(\v0/z3/z2/q2 [0]),
    .C(\v0/z3/z2/_07_ ),
    .X(\v0/z3/z2/z6/_01_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z3/z2/z6/_22_  (.A(\v0/z3/z2/_06_ ),
    .B(\v0/z3/z2/q2 [1]),
    .Y(\v0/z3/z2/z6/_02_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z3/z2/z6/_23_  (.A(\v0/z3/z2/z6/_01_ ),
    .B(\v0/z3/z2/z6/_02_ ),
    .Y(\v0/z3/z2/q5 [1]));
 sky130_fd_sc_hd__maj3_1 \v0/z3/z2/z6/_24_  (.A(\v0/z3/z2/_06_ ),
    .B(\v0/z3/z2/q2 [1]),
    .C(\v0/z3/z2/z6/_01_ ),
    .X(\v0/z3/z2/z6/_03_ ));
 sky130_fd_sc_hd__lpflow_inputiso1p_1 \v0/z3/z2/z6/_25_  (.A(\v0/z3/z2/q3 [0]),
    .SLEEP(\v0/z3/z2/q2 [2]),
    .X(\v0/z3/z2/z6/_04_ ));
 sky130_fd_sc_hd__and2_0 \v0/z3/z2/z6/_26_  (.A(\v0/z3/z2/q3 [0]),
    .B(\v0/z3/z2/q2 [2]),
    .X(\v0/z3/z2/z6/_05_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z3/z2/z6/_27_  (.A(\v0/z3/z2/q3 [0]),
    .B(\v0/z3/z2/q2 [2]),
    .Y(\v0/z3/z2/z6/_06_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z3/z2/z6/_28_  (.A(\v0/z3/z2/z6/_04_ ),
    .B(\v0/z3/z2/z6/_06_ ),
    .Y(\v0/z3/z2/z6/_07_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z3/z2/z6/_29_  (.A(\v0/z3/z2/z6/_03_ ),
    .B(\v0/z3/z2/z6/_07_ ),
    .Y(\v0/z3/z2/q5 [2]));
 sky130_fd_sc_hd__nand2_1 \v0/z3/z2/z6/_30_  (.A(\v0/z3/z2/q3 [1]),
    .B(\v0/z3/z2/q2 [3]),
    .Y(\v0/z3/z2/z6/_08_ ));
 sky130_fd_sc_hd__xor2_1 \v0/z3/z2/z6/_31_  (.A(\v0/z3/z2/q3 [1]),
    .B(\v0/z3/z2/q2 [3]),
    .X(\v0/z3/z2/z6/_09_ ));
 sky130_fd_sc_hd__o21ai_0 \v0/z3/z2/z6/_32_  (.A1(\v0/z3/z2/z6/_03_ ),
    .A2(\v0/z3/z2/z6/_05_ ),
    .B1(\v0/z3/z2/z6/_04_ ),
    .Y(\v0/z3/z2/z6/_10_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z3/z2/z6/_33_  (.A(\v0/z3/z2/z6/_09_ ),
    .B(\v0/z3/z2/z6/_10_ ),
    .Y(\v0/z3/z2/q5 [3]));
 sky130_fd_sc_hd__nor2_1 \v0/z3/z2/z6/_34_  (.A(\v0/z3/z2/q3 [2]),
    .B(\v0/z3/z2/_03_ ),
    .Y(\v0/z3/z2/z6/_11_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z3/z2/z6/_35_  (.A(\v0/z3/z2/q3 [2]),
    .B(\v0/z3/z2/_03_ ),
    .Y(\v0/z3/z2/z6/_12_ ));
 sky130_fd_sc_hd__nand2b_1 \v0/z3/z2/z6/_36_  (.A_N(\v0/z3/z2/z6/_11_ ),
    .B(\v0/z3/z2/z6/_12_ ),
    .Y(\v0/z3/z2/z6/_13_ ));
 sky130_fd_sc_hd__o221ai_1 \v0/z3/z2/z6/_37_  (.A1(\v0/z3/z2/q3 [1]),
    .A2(\v0/z3/z2/q2 [3]),
    .B1(\v0/z3/z2/z6/_03_ ),
    .B2(\v0/z3/z2/z6/_05_ ),
    .C1(\v0/z3/z2/z6/_04_ ),
    .Y(\v0/z3/z2/z6/_14_ ));
 sky130_fd_sc_hd__a21oi_1 \v0/z3/z2/z6/_38_  (.A1(\v0/z3/z2/z6/_08_ ),
    .A2(\v0/z3/z2/z6/_14_ ),
    .B1(\v0/z3/z2/z6/_13_ ),
    .Y(\v0/z3/z2/z6/_15_ ));
 sky130_fd_sc_hd__and3_1 \v0/z3/z2/z6/_39_  (.A(\v0/z3/z2/z6/_08_ ),
    .B(\v0/z3/z2/z6/_13_ ),
    .C(\v0/z3/z2/z6/_14_ ),
    .X(\v0/z3/z2/z6/_16_ ));
 sky130_fd_sc_hd__nor2_1 \v0/z3/z2/z6/_40_  (.A(\v0/z3/z2/z6/_15_ ),
    .B(\v0/z3/z2/z6/_16_ ),
    .Y(\v0/z3/z2/q5 [4]));
 sky130_fd_sc_hd__xnor2_1 \v0/z3/z2/z6/_41_  (.A(\v0/z3/z2/q3 [3]),
    .B(\v0/z3/z2/_04_ ),
    .Y(\v0/z3/z2/z6/_17_ ));
 sky130_fd_sc_hd__a31oi_1 \v0/z3/z2/z6/_42_  (.A1(\v0/z3/z2/z6/_08_ ),
    .A2(\v0/z3/z2/z6/_12_ ),
    .A3(\v0/z3/z2/z6/_14_ ),
    .B1(\v0/z3/z2/z6/_11_ ),
    .Y(\v0/z3/z2/z6/_18_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z3/z2/z6/_43_  (.A(\v0/z3/z2/z6/_17_ ),
    .B(\v0/z3/z2/z6/_18_ ),
    .Y(\v0/z3/z2/q5 [5]));
 sky130_fd_sc_hd__maj3_1 \v0/z3/z2/z6/_44_  (.A(\v0/z3/z2/q3 [3]),
    .B(\v0/z3/z2/_04_ ),
    .C(\v0/z3/z2/z6/_18_ ),
    .X(\v0/z3/z2/z6/Cout ));
 sky130_fd_sc_hd__xnor2_1 \v0/z3/z2/z7/_19_  (.A(\v0/z3/z2/q5 [0]),
    .B(\v0/z3/z2/q4 [0]),
    .Y(\v0/z3/z2/z7/_00_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z3/z2/z7/_20_  (.A(\v0/z3/z2/_10_ ),
    .B(\v0/z3/z2/z7/_00_ ),
    .Y(\v0/z3/q1 [2]));
 sky130_fd_sc_hd__maj3_1 \v0/z3/z2/z7/_21_  (.A(\v0/z3/z2/q5 [0]),
    .B(\v0/z3/z2/q4 [0]),
    .C(\v0/z3/z2/_10_ ),
    .X(\v0/z3/z2/z7/_01_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z3/z2/z7/_22_  (.A(\v0/z3/z2/q5 [1]),
    .B(\v0/z3/z2/q4 [1]),
    .Y(\v0/z3/z2/z7/_02_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z3/z2/z7/_23_  (.A(\v0/z3/z2/z7/_01_ ),
    .B(\v0/z3/z2/z7/_02_ ),
    .Y(\v0/z3/q1 [3]));
 sky130_fd_sc_hd__maj3_1 \v0/z3/z2/z7/_24_  (.A(\v0/z3/z2/q5 [1]),
    .B(\v0/z3/z2/q4 [1]),
    .C(\v0/z3/z2/z7/_01_ ),
    .X(\v0/z3/z2/z7/_03_ ));
 sky130_fd_sc_hd__lpflow_inputiso1p_1 \v0/z3/z2/z7/_25_  (.A(\v0/z3/z2/q5 [2]),
    .SLEEP(\v0/z3/z2/q4 [2]),
    .X(\v0/z3/z2/z7/_04_ ));
 sky130_fd_sc_hd__and2_0 \v0/z3/z2/z7/_26_  (.A(\v0/z3/z2/q5 [2]),
    .B(\v0/z3/z2/q4 [2]),
    .X(\v0/z3/z2/z7/_05_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z3/z2/z7/_27_  (.A(\v0/z3/z2/q5 [2]),
    .B(\v0/z3/z2/q4 [2]),
    .Y(\v0/z3/z2/z7/_06_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z3/z2/z7/_28_  (.A(\v0/z3/z2/z7/_04_ ),
    .B(\v0/z3/z2/z7/_06_ ),
    .Y(\v0/z3/z2/z7/_07_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z3/z2/z7/_29_  (.A(\v0/z3/z2/z7/_03_ ),
    .B(\v0/z3/z2/z7/_07_ ),
    .Y(\v0/z3/q1 [4]));
 sky130_fd_sc_hd__nand2_1 \v0/z3/z2/z7/_30_  (.A(\v0/z3/z2/q5 [3]),
    .B(\v0/z3/z2/q4 [3]),
    .Y(\v0/z3/z2/z7/_08_ ));
 sky130_fd_sc_hd__xor2_1 \v0/z3/z2/z7/_31_  (.A(\v0/z3/z2/q5 [3]),
    .B(\v0/z3/z2/q4 [3]),
    .X(\v0/z3/z2/z7/_09_ ));
 sky130_fd_sc_hd__o21ai_0 \v0/z3/z2/z7/_32_  (.A1(\v0/z3/z2/z7/_03_ ),
    .A2(\v0/z3/z2/z7/_05_ ),
    .B1(\v0/z3/z2/z7/_04_ ),
    .Y(\v0/z3/z2/z7/_10_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z3/z2/z7/_33_  (.A(\v0/z3/z2/z7/_09_ ),
    .B(\v0/z3/z2/z7/_10_ ),
    .Y(\v0/z3/q1 [5]));
 sky130_fd_sc_hd__nor2_1 \v0/z3/z2/z7/_34_  (.A(\v0/z3/z2/q5 [4]),
    .B(\v0/z3/z2/_08_ ),
    .Y(\v0/z3/z2/z7/_11_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z3/z2/z7/_35_  (.A(\v0/z3/z2/q5 [4]),
    .B(\v0/z3/z2/_08_ ),
    .Y(\v0/z3/z2/z7/_12_ ));
 sky130_fd_sc_hd__nand2b_1 \v0/z3/z2/z7/_36_  (.A_N(\v0/z3/z2/z7/_11_ ),
    .B(\v0/z3/z2/z7/_12_ ),
    .Y(\v0/z3/z2/z7/_13_ ));
 sky130_fd_sc_hd__o221ai_1 \v0/z3/z2/z7/_37_  (.A1(\v0/z3/z2/q5 [3]),
    .A2(\v0/z3/z2/q4 [3]),
    .B1(\v0/z3/z2/z7/_03_ ),
    .B2(\v0/z3/z2/z7/_05_ ),
    .C1(\v0/z3/z2/z7/_04_ ),
    .Y(\v0/z3/z2/z7/_14_ ));
 sky130_fd_sc_hd__a21oi_1 \v0/z3/z2/z7/_38_  (.A1(\v0/z3/z2/z7/_08_ ),
    .A2(\v0/z3/z2/z7/_14_ ),
    .B1(\v0/z3/z2/z7/_13_ ),
    .Y(\v0/z3/z2/z7/_15_ ));
 sky130_fd_sc_hd__and3_1 \v0/z3/z2/z7/_39_  (.A(\v0/z3/z2/z7/_08_ ),
    .B(\v0/z3/z2/z7/_13_ ),
    .C(\v0/z3/z2/z7/_14_ ),
    .X(\v0/z3/z2/z7/_16_ ));
 sky130_fd_sc_hd__nor2_1 \v0/z3/z2/z7/_40_  (.A(\v0/z3/z2/z7/_15_ ),
    .B(\v0/z3/z2/z7/_16_ ),
    .Y(\v0/z3/q1 [6]));
 sky130_fd_sc_hd__xnor2_1 \v0/z3/z2/z7/_41_  (.A(\v0/z3/z2/q5 [5]),
    .B(\v0/z3/z2/_09_ ),
    .Y(\v0/z3/z2/z7/_17_ ));
 sky130_fd_sc_hd__a31oi_1 \v0/z3/z2/z7/_42_  (.A1(\v0/z3/z2/z7/_08_ ),
    .A2(\v0/z3/z2/z7/_12_ ),
    .A3(\v0/z3/z2/z7/_14_ ),
    .B1(\v0/z3/z2/z7/_11_ ),
    .Y(\v0/z3/z2/z7/_18_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z3/z2/z7/_43_  (.A(\v0/z3/z2/z7/_17_ ),
    .B(\v0/z3/z2/z7/_18_ ),
    .Y(\v0/z3/q1 [7]));
 sky130_fd_sc_hd__maj3_1 \v0/z3/z2/z7/_44_  (.A(\v0/z3/z2/q5 [5]),
    .B(\v0/z3/z2/_09_ ),
    .C(\v0/z3/z2/z7/_18_ ),
    .X(\v0/z3/z2/z7/Cout ));
 sky130_fd_sc_hd__conb_1 \v0/z3/z3/_11_  (.LO(\v0/z3/z3/_00_ ));
 sky130_fd_sc_hd__conb_1 \v0/z3/z3/_12_  (.LO(\v0/z3/z3/_01_ ));
 sky130_fd_sc_hd__conb_1 \v0/z3/z3/_13_  (.LO(\v0/z3/z3/_02_ ));
 sky130_fd_sc_hd__conb_1 \v0/z3/z3/_14_  (.LO(\v0/z3/z3/_03_ ));
 sky130_fd_sc_hd__conb_1 \v0/z3/z3/_15_  (.LO(\v0/z3/z3/_04_ ));
 sky130_fd_sc_hd__conb_1 \v0/z3/z3/_16_  (.LO(\v0/z3/z3/_05_ ));
 sky130_fd_sc_hd__conb_1 \v0/z3/z3/_17_  (.LO(\v0/z3/z3/_06_ ));
 sky130_fd_sc_hd__conb_1 \v0/z3/z3/_18_  (.LO(\v0/z3/z3/_07_ ));
 sky130_fd_sc_hd__conb_1 \v0/z3/z3/_19_  (.LO(\v0/z3/z3/_08_ ));
 sky130_fd_sc_hd__conb_1 \v0/z3/z3/_20_  (.LO(\v0/z3/z3/_09_ ));
 sky130_fd_sc_hd__conb_1 \v0/z3/z3/_21_  (.LO(\v0/z3/z3/_10_ ));
 sky130_fd_sc_hd__and2_0 \v0/z3/z3/z1/_0_  (.A(abs_b[12]),
    .B(a[0]),
    .X(\v0/z3/q2 [0]));
 sky130_fd_sc_hd__and2_0 \v0/z3/z3/z1/_1_  (.A(abs_b[12]),
    .B(abs_a[1]),
    .X(\v0/z3/z3/z1/temp [0]));
 sky130_fd_sc_hd__and2_0 \v0/z3/z3/z1/_2_  (.A(a[0]),
    .B(abs_b[13]),
    .X(\v0/z3/z3/z1/temp [1]));
 sky130_fd_sc_hd__and2_0 \v0/z3/z3/z1/_3_  (.A(abs_a[1]),
    .B(abs_b[13]),
    .X(\v0/z3/z3/z1/temp [2]));
 sky130_fd_sc_hd__and2_0 \v0/z3/z3/z1/z1/_0_  (.A(\v0/z3/z3/z1/temp [1]),
    .B(\v0/z3/z3/z1/temp [0]),
    .X(\v0/z3/z3/z1/temp [3]));
 sky130_fd_sc_hd__xor2_1 \v0/z3/z3/z1/z1/_1_  (.A(\v0/z3/z3/z1/temp [1]),
    .B(\v0/z3/z3/z1/temp [0]),
    .X(\v0/z3/q2 [1]));
 sky130_fd_sc_hd__and2_0 \v0/z3/z3/z1/z2/_0_  (.A(\v0/z3/z3/z1/temp [3]),
    .B(\v0/z3/z3/z1/temp [2]),
    .X(\v0/z3/z3/q0 [3]));
 sky130_fd_sc_hd__xor2_1 \v0/z3/z3/z1/z2/_1_  (.A(\v0/z3/z3/z1/temp [3]),
    .B(\v0/z3/z3/z1/temp [2]),
    .X(\v0/z3/z3/q0 [2]));
 sky130_fd_sc_hd__and2_0 \v0/z3/z3/z2/_0_  (.A(abs_b[12]),
    .B(abs_a[2]),
    .X(\v0/z3/z3/q1 [0]));
 sky130_fd_sc_hd__and2_0 \v0/z3/z3/z2/_1_  (.A(abs_b[12]),
    .B(abs_a[3]),
    .X(\v0/z3/z3/z2/temp [0]));
 sky130_fd_sc_hd__and2_0 \v0/z3/z3/z2/_2_  (.A(abs_a[2]),
    .B(abs_b[13]),
    .X(\v0/z3/z3/z2/temp [1]));
 sky130_fd_sc_hd__and2_0 \v0/z3/z3/z2/_3_  (.A(abs_a[3]),
    .B(abs_b[13]),
    .X(\v0/z3/z3/z2/temp [2]));
 sky130_fd_sc_hd__and2_0 \v0/z3/z3/z2/z1/_0_  (.A(\v0/z3/z3/z2/temp [1]),
    .B(\v0/z3/z3/z2/temp [0]),
    .X(\v0/z3/z3/z2/temp [3]));
 sky130_fd_sc_hd__xor2_1 \v0/z3/z3/z2/z1/_1_  (.A(\v0/z3/z3/z2/temp [1]),
    .B(\v0/z3/z3/z2/temp [0]),
    .X(\v0/z3/z3/q1 [1]));
 sky130_fd_sc_hd__and2_0 \v0/z3/z3/z2/z2/_0_  (.A(\v0/z3/z3/z2/temp [3]),
    .B(\v0/z3/z3/z2/temp [2]),
    .X(\v0/z3/z3/q1 [3]));
 sky130_fd_sc_hd__xor2_1 \v0/z3/z3/z2/z2/_1_  (.A(\v0/z3/z3/z2/temp [3]),
    .B(\v0/z3/z3/z2/temp [2]),
    .X(\v0/z3/z3/q1 [2]));
 sky130_fd_sc_hd__and2_0 \v0/z3/z3/z3/_0_  (.A(abs_b[14]),
    .B(a[0]),
    .X(\v0/z3/z3/q2 [0]));
 sky130_fd_sc_hd__and2_0 \v0/z3/z3/z3/_1_  (.A(abs_b[14]),
    .B(abs_a[1]),
    .X(\v0/z3/z3/z3/temp [0]));
 sky130_fd_sc_hd__and2_0 \v0/z3/z3/z3/_2_  (.A(a[0]),
    .B(abs_b[15]),
    .X(\v0/z3/z3/z3/temp [1]));
 sky130_fd_sc_hd__and2_0 \v0/z3/z3/z3/_3_  (.A(abs_a[1]),
    .B(abs_b[15]),
    .X(\v0/z3/z3/z3/temp [2]));
 sky130_fd_sc_hd__and2_0 \v0/z3/z3/z3/z1/_0_  (.A(\v0/z3/z3/z3/temp [1]),
    .B(\v0/z3/z3/z3/temp [0]),
    .X(\v0/z3/z3/z3/temp [3]));
 sky130_fd_sc_hd__xor2_1 \v0/z3/z3/z3/z1/_1_  (.A(\v0/z3/z3/z3/temp [1]),
    .B(\v0/z3/z3/z3/temp [0]),
    .X(\v0/z3/z3/q2 [1]));
 sky130_fd_sc_hd__and2_0 \v0/z3/z3/z3/z2/_0_  (.A(\v0/z3/z3/z3/temp [3]),
    .B(\v0/z3/z3/z3/temp [2]),
    .X(\v0/z3/z3/q2 [3]));
 sky130_fd_sc_hd__xor2_1 \v0/z3/z3/z3/z2/_1_  (.A(\v0/z3/z3/z3/temp [3]),
    .B(\v0/z3/z3/z3/temp [2]),
    .X(\v0/z3/z3/q2 [2]));
 sky130_fd_sc_hd__and2_0 \v0/z3/z3/z4/_0_  (.A(abs_b[14]),
    .B(abs_a[2]),
    .X(\v0/z3/z3/q3 [0]));
 sky130_fd_sc_hd__and2_0 \v0/z3/z3/z4/_1_  (.A(abs_b[14]),
    .B(abs_a[3]),
    .X(\v0/z3/z3/z4/temp [0]));
 sky130_fd_sc_hd__and2_0 \v0/z3/z3/z4/_2_  (.A(abs_a[2]),
    .B(abs_b[15]),
    .X(\v0/z3/z3/z4/temp [1]));
 sky130_fd_sc_hd__and2_0 \v0/z3/z3/z4/_3_  (.A(abs_a[3]),
    .B(abs_b[15]),
    .X(\v0/z3/z3/z4/temp [2]));
 sky130_fd_sc_hd__and2_0 \v0/z3/z3/z4/z1/_0_  (.A(\v0/z3/z3/z4/temp [1]),
    .B(\v0/z3/z3/z4/temp [0]),
    .X(\v0/z3/z3/z4/temp [3]));
 sky130_fd_sc_hd__xor2_1 \v0/z3/z3/z4/z1/_1_  (.A(\v0/z3/z3/z4/temp [1]),
    .B(\v0/z3/z3/z4/temp [0]),
    .X(\v0/z3/z3/q3 [1]));
 sky130_fd_sc_hd__and2_0 \v0/z3/z3/z4/z2/_0_  (.A(\v0/z3/z3/z4/temp [3]),
    .B(\v0/z3/z3/z4/temp [2]),
    .X(\v0/z3/z3/q3 [3]));
 sky130_fd_sc_hd__xor2_1 \v0/z3/z3/z4/z2/_1_  (.A(\v0/z3/z3/z4/temp [3]),
    .B(\v0/z3/z3/z4/temp [2]),
    .X(\v0/z3/z3/q3 [2]));
 sky130_fd_sc_hd__xnor2_1 \v0/z3/z3/z5/_07_  (.A(\v0/z3/z3/q0 [2]),
    .B(\v0/z3/z3/q1 [0]),
    .Y(\v0/z3/z3/z5/_00_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z3/z3/z5/_08_  (.A(\v0/z3/z3/_02_ ),
    .B(\v0/z3/z3/z5/_00_ ),
    .Y(\v0/z3/z3/q4 [0]));
 sky130_fd_sc_hd__maj3_1 \v0/z3/z3/z5/_09_  (.A(\v0/z3/z3/q0 [2]),
    .B(\v0/z3/z3/q1 [0]),
    .C(\v0/z3/z3/_02_ ),
    .X(\v0/z3/z3/z5/_01_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z3/z3/z5/_10_  (.A(\v0/z3/z3/q0 [3]),
    .B(\v0/z3/z3/q1 [1]),
    .Y(\v0/z3/z3/z5/_02_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z3/z3/z5/_11_  (.A(\v0/z3/z3/z5/_01_ ),
    .B(\v0/z3/z3/z5/_02_ ),
    .Y(\v0/z3/z3/q4 [1]));
 sky130_fd_sc_hd__maj3_1 \v0/z3/z3/z5/_12_  (.A(\v0/z3/z3/q0 [3]),
    .B(\v0/z3/z3/q1 [1]),
    .C(\v0/z3/z3/z5/_01_ ),
    .X(\v0/z3/z3/z5/_03_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z3/z3/z5/_13_  (.A(\v0/z3/z3/_00_ ),
    .B(\v0/z3/z3/q1 [2]),
    .Y(\v0/z3/z3/z5/_04_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z3/z3/z5/_14_  (.A(\v0/z3/z3/z5/_03_ ),
    .B(\v0/z3/z3/z5/_04_ ),
    .Y(\v0/z3/z3/q4 [2]));
 sky130_fd_sc_hd__maj3_1 \v0/z3/z3/z5/_15_  (.A(\v0/z3/z3/_00_ ),
    .B(\v0/z3/z3/q1 [2]),
    .C(\v0/z3/z3/z5/_03_ ),
    .X(\v0/z3/z3/z5/_05_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z3/z3/z5/_16_  (.A(\v0/z3/z3/_01_ ),
    .B(\v0/z3/z3/q1 [3]),
    .Y(\v0/z3/z3/z5/_06_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z3/z3/z5/_17_  (.A(\v0/z3/z3/z5/_05_ ),
    .B(\v0/z3/z3/z5/_06_ ),
    .Y(\v0/z3/z3/q4 [3]));
 sky130_fd_sc_hd__maj3_1 \v0/z3/z3/z5/_18_  (.A(\v0/z3/z3/_01_ ),
    .B(\v0/z3/z3/q1 [3]),
    .C(\v0/z3/z3/z5/_05_ ),
    .X(\v0/z3/z3/z5/Cout ));
 sky130_fd_sc_hd__xnor2_1 \v0/z3/z3/z6/_19_  (.A(\v0/z3/z3/_05_ ),
    .B(\v0/z3/z3/q2 [0]),
    .Y(\v0/z3/z3/z6/_00_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z3/z3/z6/_20_  (.A(\v0/z3/z3/_07_ ),
    .B(\v0/z3/z3/z6/_00_ ),
    .Y(\v0/z3/z3/q5 [0]));
 sky130_fd_sc_hd__maj3_1 \v0/z3/z3/z6/_21_  (.A(\v0/z3/z3/_05_ ),
    .B(\v0/z3/z3/q2 [0]),
    .C(\v0/z3/z3/_07_ ),
    .X(\v0/z3/z3/z6/_01_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z3/z3/z6/_22_  (.A(\v0/z3/z3/_06_ ),
    .B(\v0/z3/z3/q2 [1]),
    .Y(\v0/z3/z3/z6/_02_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z3/z3/z6/_23_  (.A(\v0/z3/z3/z6/_01_ ),
    .B(\v0/z3/z3/z6/_02_ ),
    .Y(\v0/z3/z3/q5 [1]));
 sky130_fd_sc_hd__maj3_1 \v0/z3/z3/z6/_24_  (.A(\v0/z3/z3/_06_ ),
    .B(\v0/z3/z3/q2 [1]),
    .C(\v0/z3/z3/z6/_01_ ),
    .X(\v0/z3/z3/z6/_03_ ));
 sky130_fd_sc_hd__lpflow_inputiso1p_1 \v0/z3/z3/z6/_25_  (.A(\v0/z3/z3/q3 [0]),
    .SLEEP(\v0/z3/z3/q2 [2]),
    .X(\v0/z3/z3/z6/_04_ ));
 sky130_fd_sc_hd__and2_0 \v0/z3/z3/z6/_26_  (.A(\v0/z3/z3/q3 [0]),
    .B(\v0/z3/z3/q2 [2]),
    .X(\v0/z3/z3/z6/_05_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z3/z3/z6/_27_  (.A(\v0/z3/z3/q3 [0]),
    .B(\v0/z3/z3/q2 [2]),
    .Y(\v0/z3/z3/z6/_06_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z3/z3/z6/_28_  (.A(\v0/z3/z3/z6/_04_ ),
    .B(\v0/z3/z3/z6/_06_ ),
    .Y(\v0/z3/z3/z6/_07_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z3/z3/z6/_29_  (.A(\v0/z3/z3/z6/_03_ ),
    .B(\v0/z3/z3/z6/_07_ ),
    .Y(\v0/z3/z3/q5 [2]));
 sky130_fd_sc_hd__nand2_1 \v0/z3/z3/z6/_30_  (.A(\v0/z3/z3/q3 [1]),
    .B(\v0/z3/z3/q2 [3]),
    .Y(\v0/z3/z3/z6/_08_ ));
 sky130_fd_sc_hd__xor2_1 \v0/z3/z3/z6/_31_  (.A(\v0/z3/z3/q3 [1]),
    .B(\v0/z3/z3/q2 [3]),
    .X(\v0/z3/z3/z6/_09_ ));
 sky130_fd_sc_hd__o21ai_0 \v0/z3/z3/z6/_32_  (.A1(\v0/z3/z3/z6/_03_ ),
    .A2(\v0/z3/z3/z6/_05_ ),
    .B1(\v0/z3/z3/z6/_04_ ),
    .Y(\v0/z3/z3/z6/_10_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z3/z3/z6/_33_  (.A(\v0/z3/z3/z6/_09_ ),
    .B(\v0/z3/z3/z6/_10_ ),
    .Y(\v0/z3/z3/q5 [3]));
 sky130_fd_sc_hd__nor2_1 \v0/z3/z3/z6/_34_  (.A(\v0/z3/z3/q3 [2]),
    .B(\v0/z3/z3/_03_ ),
    .Y(\v0/z3/z3/z6/_11_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z3/z3/z6/_35_  (.A(\v0/z3/z3/q3 [2]),
    .B(\v0/z3/z3/_03_ ),
    .Y(\v0/z3/z3/z6/_12_ ));
 sky130_fd_sc_hd__nand2b_1 \v0/z3/z3/z6/_36_  (.A_N(\v0/z3/z3/z6/_11_ ),
    .B(\v0/z3/z3/z6/_12_ ),
    .Y(\v0/z3/z3/z6/_13_ ));
 sky130_fd_sc_hd__o221ai_1 \v0/z3/z3/z6/_37_  (.A1(\v0/z3/z3/q3 [1]),
    .A2(\v0/z3/z3/q2 [3]),
    .B1(\v0/z3/z3/z6/_03_ ),
    .B2(\v0/z3/z3/z6/_05_ ),
    .C1(\v0/z3/z3/z6/_04_ ),
    .Y(\v0/z3/z3/z6/_14_ ));
 sky130_fd_sc_hd__a21oi_1 \v0/z3/z3/z6/_38_  (.A1(\v0/z3/z3/z6/_08_ ),
    .A2(\v0/z3/z3/z6/_14_ ),
    .B1(\v0/z3/z3/z6/_13_ ),
    .Y(\v0/z3/z3/z6/_15_ ));
 sky130_fd_sc_hd__and3_1 \v0/z3/z3/z6/_39_  (.A(\v0/z3/z3/z6/_08_ ),
    .B(\v0/z3/z3/z6/_13_ ),
    .C(\v0/z3/z3/z6/_14_ ),
    .X(\v0/z3/z3/z6/_16_ ));
 sky130_fd_sc_hd__nor2_1 \v0/z3/z3/z6/_40_  (.A(\v0/z3/z3/z6/_15_ ),
    .B(\v0/z3/z3/z6/_16_ ),
    .Y(\v0/z3/z3/q5 [4]));
 sky130_fd_sc_hd__xnor2_1 \v0/z3/z3/z6/_41_  (.A(\v0/z3/z3/q3 [3]),
    .B(\v0/z3/z3/_04_ ),
    .Y(\v0/z3/z3/z6/_17_ ));
 sky130_fd_sc_hd__a31oi_1 \v0/z3/z3/z6/_42_  (.A1(\v0/z3/z3/z6/_08_ ),
    .A2(\v0/z3/z3/z6/_12_ ),
    .A3(\v0/z3/z3/z6/_14_ ),
    .B1(\v0/z3/z3/z6/_11_ ),
    .Y(\v0/z3/z3/z6/_18_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z3/z3/z6/_43_  (.A(\v0/z3/z3/z6/_17_ ),
    .B(\v0/z3/z3/z6/_18_ ),
    .Y(\v0/z3/z3/q5 [5]));
 sky130_fd_sc_hd__maj3_1 \v0/z3/z3/z6/_44_  (.A(\v0/z3/z3/q3 [3]),
    .B(\v0/z3/z3/_04_ ),
    .C(\v0/z3/z3/z6/_18_ ),
    .X(\v0/z3/z3/z6/Cout ));
 sky130_fd_sc_hd__xnor2_1 \v0/z3/z3/z7/_19_  (.A(\v0/z3/z3/q5 [0]),
    .B(\v0/z3/z3/q4 [0]),
    .Y(\v0/z3/z3/z7/_00_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z3/z3/z7/_20_  (.A(\v0/z3/z3/_10_ ),
    .B(\v0/z3/z3/z7/_00_ ),
    .Y(\v0/z3/q2 [2]));
 sky130_fd_sc_hd__maj3_1 \v0/z3/z3/z7/_21_  (.A(\v0/z3/z3/q5 [0]),
    .B(\v0/z3/z3/q4 [0]),
    .C(\v0/z3/z3/_10_ ),
    .X(\v0/z3/z3/z7/_01_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z3/z3/z7/_22_  (.A(\v0/z3/z3/q5 [1]),
    .B(\v0/z3/z3/q4 [1]),
    .Y(\v0/z3/z3/z7/_02_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z3/z3/z7/_23_  (.A(\v0/z3/z3/z7/_01_ ),
    .B(\v0/z3/z3/z7/_02_ ),
    .Y(\v0/z3/q2 [3]));
 sky130_fd_sc_hd__maj3_1 \v0/z3/z3/z7/_24_  (.A(\v0/z3/z3/q5 [1]),
    .B(\v0/z3/z3/q4 [1]),
    .C(\v0/z3/z3/z7/_01_ ),
    .X(\v0/z3/z3/z7/_03_ ));
 sky130_fd_sc_hd__lpflow_inputiso1p_1 \v0/z3/z3/z7/_25_  (.A(\v0/z3/z3/q5 [2]),
    .SLEEP(\v0/z3/z3/q4 [2]),
    .X(\v0/z3/z3/z7/_04_ ));
 sky130_fd_sc_hd__and2_0 \v0/z3/z3/z7/_26_  (.A(\v0/z3/z3/q5 [2]),
    .B(\v0/z3/z3/q4 [2]),
    .X(\v0/z3/z3/z7/_05_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z3/z3/z7/_27_  (.A(\v0/z3/z3/q5 [2]),
    .B(\v0/z3/z3/q4 [2]),
    .Y(\v0/z3/z3/z7/_06_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z3/z3/z7/_28_  (.A(\v0/z3/z3/z7/_04_ ),
    .B(\v0/z3/z3/z7/_06_ ),
    .Y(\v0/z3/z3/z7/_07_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z3/z3/z7/_29_  (.A(\v0/z3/z3/z7/_03_ ),
    .B(\v0/z3/z3/z7/_07_ ),
    .Y(\v0/z3/q2 [4]));
 sky130_fd_sc_hd__nand2_1 \v0/z3/z3/z7/_30_  (.A(\v0/z3/z3/q5 [3]),
    .B(\v0/z3/z3/q4 [3]),
    .Y(\v0/z3/z3/z7/_08_ ));
 sky130_fd_sc_hd__xor2_1 \v0/z3/z3/z7/_31_  (.A(\v0/z3/z3/q5 [3]),
    .B(\v0/z3/z3/q4 [3]),
    .X(\v0/z3/z3/z7/_09_ ));
 sky130_fd_sc_hd__o21ai_0 \v0/z3/z3/z7/_32_  (.A1(\v0/z3/z3/z7/_03_ ),
    .A2(\v0/z3/z3/z7/_05_ ),
    .B1(\v0/z3/z3/z7/_04_ ),
    .Y(\v0/z3/z3/z7/_10_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z3/z3/z7/_33_  (.A(\v0/z3/z3/z7/_09_ ),
    .B(\v0/z3/z3/z7/_10_ ),
    .Y(\v0/z3/q2 [5]));
 sky130_fd_sc_hd__nor2_1 \v0/z3/z3/z7/_34_  (.A(\v0/z3/z3/q5 [4]),
    .B(\v0/z3/z3/_08_ ),
    .Y(\v0/z3/z3/z7/_11_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z3/z3/z7/_35_  (.A(\v0/z3/z3/q5 [4]),
    .B(\v0/z3/z3/_08_ ),
    .Y(\v0/z3/z3/z7/_12_ ));
 sky130_fd_sc_hd__nand2b_1 \v0/z3/z3/z7/_36_  (.A_N(\v0/z3/z3/z7/_11_ ),
    .B(\v0/z3/z3/z7/_12_ ),
    .Y(\v0/z3/z3/z7/_13_ ));
 sky130_fd_sc_hd__o221ai_1 \v0/z3/z3/z7/_37_  (.A1(\v0/z3/z3/q5 [3]),
    .A2(\v0/z3/z3/q4 [3]),
    .B1(\v0/z3/z3/z7/_03_ ),
    .B2(\v0/z3/z3/z7/_05_ ),
    .C1(\v0/z3/z3/z7/_04_ ),
    .Y(\v0/z3/z3/z7/_14_ ));
 sky130_fd_sc_hd__a21oi_1 \v0/z3/z3/z7/_38_  (.A1(\v0/z3/z3/z7/_08_ ),
    .A2(\v0/z3/z3/z7/_14_ ),
    .B1(\v0/z3/z3/z7/_13_ ),
    .Y(\v0/z3/z3/z7/_15_ ));
 sky130_fd_sc_hd__and3_1 \v0/z3/z3/z7/_39_  (.A(\v0/z3/z3/z7/_08_ ),
    .B(\v0/z3/z3/z7/_13_ ),
    .C(\v0/z3/z3/z7/_14_ ),
    .X(\v0/z3/z3/z7/_16_ ));
 sky130_fd_sc_hd__nor2_1 \v0/z3/z3/z7/_40_  (.A(\v0/z3/z3/z7/_15_ ),
    .B(\v0/z3/z3/z7/_16_ ),
    .Y(\v0/z3/q2 [6]));
 sky130_fd_sc_hd__xnor2_1 \v0/z3/z3/z7/_41_  (.A(\v0/z3/z3/q5 [5]),
    .B(\v0/z3/z3/_09_ ),
    .Y(\v0/z3/z3/z7/_17_ ));
 sky130_fd_sc_hd__a31oi_1 \v0/z3/z3/z7/_42_  (.A1(\v0/z3/z3/z7/_08_ ),
    .A2(\v0/z3/z3/z7/_12_ ),
    .A3(\v0/z3/z3/z7/_14_ ),
    .B1(\v0/z3/z3/z7/_11_ ),
    .Y(\v0/z3/z3/z7/_18_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z3/z3/z7/_43_  (.A(\v0/z3/z3/z7/_17_ ),
    .B(\v0/z3/z3/z7/_18_ ),
    .Y(\v0/z3/q2 [7]));
 sky130_fd_sc_hd__maj3_1 \v0/z3/z3/z7/_44_  (.A(\v0/z3/z3/q5 [5]),
    .B(\v0/z3/z3/_09_ ),
    .C(\v0/z3/z3/z7/_18_ ),
    .X(\v0/z3/z3/z7/Cout ));
 sky130_fd_sc_hd__conb_1 \v0/z3/z4/_11_  (.LO(\v0/z3/z4/_00_ ));
 sky130_fd_sc_hd__conb_1 \v0/z3/z4/_12_  (.LO(\v0/z3/z4/_01_ ));
 sky130_fd_sc_hd__conb_1 \v0/z3/z4/_13_  (.LO(\v0/z3/z4/_02_ ));
 sky130_fd_sc_hd__conb_1 \v0/z3/z4/_14_  (.LO(\v0/z3/z4/_03_ ));
 sky130_fd_sc_hd__conb_1 \v0/z3/z4/_15_  (.LO(\v0/z3/z4/_04_ ));
 sky130_fd_sc_hd__conb_1 \v0/z3/z4/_16_  (.LO(\v0/z3/z4/_05_ ));
 sky130_fd_sc_hd__conb_1 \v0/z3/z4/_17_  (.LO(\v0/z3/z4/_06_ ));
 sky130_fd_sc_hd__conb_1 \v0/z3/z4/_18_  (.LO(\v0/z3/z4/_07_ ));
 sky130_fd_sc_hd__conb_1 \v0/z3/z4/_19_  (.LO(\v0/z3/z4/_08_ ));
 sky130_fd_sc_hd__conb_1 \v0/z3/z4/_20_  (.LO(\v0/z3/z4/_09_ ));
 sky130_fd_sc_hd__conb_1 \v0/z3/z4/_21_  (.LO(\v0/z3/z4/_10_ ));
 sky130_fd_sc_hd__and2_0 \v0/z3/z4/z1/_0_  (.A(abs_b[12]),
    .B(abs_a[4]),
    .X(\v0/z3/q3 [0]));
 sky130_fd_sc_hd__and2_0 \v0/z3/z4/z1/_1_  (.A(abs_b[12]),
    .B(abs_a[5]),
    .X(\v0/z3/z4/z1/temp [0]));
 sky130_fd_sc_hd__and2_0 \v0/z3/z4/z1/_2_  (.A(abs_a[4]),
    .B(abs_b[13]),
    .X(\v0/z3/z4/z1/temp [1]));
 sky130_fd_sc_hd__and2_0 \v0/z3/z4/z1/_3_  (.A(abs_a[5]),
    .B(abs_b[13]),
    .X(\v0/z3/z4/z1/temp [2]));
 sky130_fd_sc_hd__and2_0 \v0/z3/z4/z1/z1/_0_  (.A(\v0/z3/z4/z1/temp [1]),
    .B(\v0/z3/z4/z1/temp [0]),
    .X(\v0/z3/z4/z1/temp [3]));
 sky130_fd_sc_hd__xor2_1 \v0/z3/z4/z1/z1/_1_  (.A(\v0/z3/z4/z1/temp [1]),
    .B(\v0/z3/z4/z1/temp [0]),
    .X(\v0/z3/q3 [1]));
 sky130_fd_sc_hd__and2_0 \v0/z3/z4/z1/z2/_0_  (.A(\v0/z3/z4/z1/temp [3]),
    .B(\v0/z3/z4/z1/temp [2]),
    .X(\v0/z3/z4/q0 [3]));
 sky130_fd_sc_hd__xor2_1 \v0/z3/z4/z1/z2/_1_  (.A(\v0/z3/z4/z1/temp [3]),
    .B(\v0/z3/z4/z1/temp [2]),
    .X(\v0/z3/z4/q0 [2]));
 sky130_fd_sc_hd__and2_0 \v0/z3/z4/z2/_0_  (.A(abs_b[12]),
    .B(abs_a[6]),
    .X(\v0/z3/z4/q1 [0]));
 sky130_fd_sc_hd__and2_0 \v0/z3/z4/z2/_1_  (.A(abs_b[12]),
    .B(abs_a[7]),
    .X(\v0/z3/z4/z2/temp [0]));
 sky130_fd_sc_hd__and2_0 \v0/z3/z4/z2/_2_  (.A(abs_a[6]),
    .B(abs_b[13]),
    .X(\v0/z3/z4/z2/temp [1]));
 sky130_fd_sc_hd__and2_0 \v0/z3/z4/z2/_3_  (.A(abs_a[7]),
    .B(abs_b[13]),
    .X(\v0/z3/z4/z2/temp [2]));
 sky130_fd_sc_hd__and2_0 \v0/z3/z4/z2/z1/_0_  (.A(\v0/z3/z4/z2/temp [1]),
    .B(\v0/z3/z4/z2/temp [0]),
    .X(\v0/z3/z4/z2/temp [3]));
 sky130_fd_sc_hd__xor2_1 \v0/z3/z4/z2/z1/_1_  (.A(\v0/z3/z4/z2/temp [1]),
    .B(\v0/z3/z4/z2/temp [0]),
    .X(\v0/z3/z4/q1 [1]));
 sky130_fd_sc_hd__and2_0 \v0/z3/z4/z2/z2/_0_  (.A(\v0/z3/z4/z2/temp [3]),
    .B(\v0/z3/z4/z2/temp [2]),
    .X(\v0/z3/z4/q1 [3]));
 sky130_fd_sc_hd__xor2_1 \v0/z3/z4/z2/z2/_1_  (.A(\v0/z3/z4/z2/temp [3]),
    .B(\v0/z3/z4/z2/temp [2]),
    .X(\v0/z3/z4/q1 [2]));
 sky130_fd_sc_hd__and2_0 \v0/z3/z4/z3/_0_  (.A(abs_b[14]),
    .B(abs_a[4]),
    .X(\v0/z3/z4/q2 [0]));
 sky130_fd_sc_hd__and2_0 \v0/z3/z4/z3/_1_  (.A(abs_b[14]),
    .B(abs_a[5]),
    .X(\v0/z3/z4/z3/temp [0]));
 sky130_fd_sc_hd__and2_0 \v0/z3/z4/z3/_2_  (.A(abs_a[4]),
    .B(abs_b[15]),
    .X(\v0/z3/z4/z3/temp [1]));
 sky130_fd_sc_hd__and2_0 \v0/z3/z4/z3/_3_  (.A(abs_a[5]),
    .B(abs_b[15]),
    .X(\v0/z3/z4/z3/temp [2]));
 sky130_fd_sc_hd__and2_0 \v0/z3/z4/z3/z1/_0_  (.A(\v0/z3/z4/z3/temp [1]),
    .B(\v0/z3/z4/z3/temp [0]),
    .X(\v0/z3/z4/z3/temp [3]));
 sky130_fd_sc_hd__xor2_1 \v0/z3/z4/z3/z1/_1_  (.A(\v0/z3/z4/z3/temp [1]),
    .B(\v0/z3/z4/z3/temp [0]),
    .X(\v0/z3/z4/q2 [1]));
 sky130_fd_sc_hd__and2_0 \v0/z3/z4/z3/z2/_0_  (.A(\v0/z3/z4/z3/temp [3]),
    .B(\v0/z3/z4/z3/temp [2]),
    .X(\v0/z3/z4/q2 [3]));
 sky130_fd_sc_hd__xor2_1 \v0/z3/z4/z3/z2/_1_  (.A(\v0/z3/z4/z3/temp [3]),
    .B(\v0/z3/z4/z3/temp [2]),
    .X(\v0/z3/z4/q2 [2]));
 sky130_fd_sc_hd__and2_0 \v0/z3/z4/z4/_0_  (.A(abs_b[14]),
    .B(abs_a[6]),
    .X(\v0/z3/z4/q3 [0]));
 sky130_fd_sc_hd__and2_0 \v0/z3/z4/z4/_1_  (.A(abs_b[14]),
    .B(abs_a[7]),
    .X(\v0/z3/z4/z4/temp [0]));
 sky130_fd_sc_hd__and2_0 \v0/z3/z4/z4/_2_  (.A(abs_a[6]),
    .B(abs_b[15]),
    .X(\v0/z3/z4/z4/temp [1]));
 sky130_fd_sc_hd__and2_0 \v0/z3/z4/z4/_3_  (.A(abs_a[7]),
    .B(abs_b[15]),
    .X(\v0/z3/z4/z4/temp [2]));
 sky130_fd_sc_hd__and2_0 \v0/z3/z4/z4/z1/_0_  (.A(\v0/z3/z4/z4/temp [1]),
    .B(\v0/z3/z4/z4/temp [0]),
    .X(\v0/z3/z4/z4/temp [3]));
 sky130_fd_sc_hd__xor2_1 \v0/z3/z4/z4/z1/_1_  (.A(\v0/z3/z4/z4/temp [1]),
    .B(\v0/z3/z4/z4/temp [0]),
    .X(\v0/z3/z4/q3 [1]));
 sky130_fd_sc_hd__and2_0 \v0/z3/z4/z4/z2/_0_  (.A(\v0/z3/z4/z4/temp [3]),
    .B(\v0/z3/z4/z4/temp [2]),
    .X(\v0/z3/z4/q3 [3]));
 sky130_fd_sc_hd__xor2_1 \v0/z3/z4/z4/z2/_1_  (.A(\v0/z3/z4/z4/temp [3]),
    .B(\v0/z3/z4/z4/temp [2]),
    .X(\v0/z3/z4/q3 [2]));
 sky130_fd_sc_hd__xnor2_1 \v0/z3/z4/z5/_07_  (.A(\v0/z3/z4/q0 [2]),
    .B(\v0/z3/z4/q1 [0]),
    .Y(\v0/z3/z4/z5/_00_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z3/z4/z5/_08_  (.A(\v0/z3/z4/_02_ ),
    .B(\v0/z3/z4/z5/_00_ ),
    .Y(\v0/z3/z4/q4 [0]));
 sky130_fd_sc_hd__maj3_1 \v0/z3/z4/z5/_09_  (.A(\v0/z3/z4/q0 [2]),
    .B(\v0/z3/z4/q1 [0]),
    .C(\v0/z3/z4/_02_ ),
    .X(\v0/z3/z4/z5/_01_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z3/z4/z5/_10_  (.A(\v0/z3/z4/q0 [3]),
    .B(\v0/z3/z4/q1 [1]),
    .Y(\v0/z3/z4/z5/_02_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z3/z4/z5/_11_  (.A(\v0/z3/z4/z5/_01_ ),
    .B(\v0/z3/z4/z5/_02_ ),
    .Y(\v0/z3/z4/q4 [1]));
 sky130_fd_sc_hd__maj3_1 \v0/z3/z4/z5/_12_  (.A(\v0/z3/z4/q0 [3]),
    .B(\v0/z3/z4/q1 [1]),
    .C(\v0/z3/z4/z5/_01_ ),
    .X(\v0/z3/z4/z5/_03_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z3/z4/z5/_13_  (.A(\v0/z3/z4/_00_ ),
    .B(\v0/z3/z4/q1 [2]),
    .Y(\v0/z3/z4/z5/_04_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z3/z4/z5/_14_  (.A(\v0/z3/z4/z5/_03_ ),
    .B(\v0/z3/z4/z5/_04_ ),
    .Y(\v0/z3/z4/q4 [2]));
 sky130_fd_sc_hd__maj3_1 \v0/z3/z4/z5/_15_  (.A(\v0/z3/z4/_00_ ),
    .B(\v0/z3/z4/q1 [2]),
    .C(\v0/z3/z4/z5/_03_ ),
    .X(\v0/z3/z4/z5/_05_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z3/z4/z5/_16_  (.A(\v0/z3/z4/_01_ ),
    .B(\v0/z3/z4/q1 [3]),
    .Y(\v0/z3/z4/z5/_06_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z3/z4/z5/_17_  (.A(\v0/z3/z4/z5/_05_ ),
    .B(\v0/z3/z4/z5/_06_ ),
    .Y(\v0/z3/z4/q4 [3]));
 sky130_fd_sc_hd__maj3_1 \v0/z3/z4/z5/_18_  (.A(\v0/z3/z4/_01_ ),
    .B(\v0/z3/z4/q1 [3]),
    .C(\v0/z3/z4/z5/_05_ ),
    .X(\v0/z3/z4/z5/Cout ));
 sky130_fd_sc_hd__xnor2_1 \v0/z3/z4/z6/_19_  (.A(\v0/z3/z4/_05_ ),
    .B(\v0/z3/z4/q2 [0]),
    .Y(\v0/z3/z4/z6/_00_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z3/z4/z6/_20_  (.A(\v0/z3/z4/_07_ ),
    .B(\v0/z3/z4/z6/_00_ ),
    .Y(\v0/z3/z4/q5 [0]));
 sky130_fd_sc_hd__maj3_1 \v0/z3/z4/z6/_21_  (.A(\v0/z3/z4/_05_ ),
    .B(\v0/z3/z4/q2 [0]),
    .C(\v0/z3/z4/_07_ ),
    .X(\v0/z3/z4/z6/_01_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z3/z4/z6/_22_  (.A(\v0/z3/z4/_06_ ),
    .B(\v0/z3/z4/q2 [1]),
    .Y(\v0/z3/z4/z6/_02_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z3/z4/z6/_23_  (.A(\v0/z3/z4/z6/_01_ ),
    .B(\v0/z3/z4/z6/_02_ ),
    .Y(\v0/z3/z4/q5 [1]));
 sky130_fd_sc_hd__maj3_1 \v0/z3/z4/z6/_24_  (.A(\v0/z3/z4/_06_ ),
    .B(\v0/z3/z4/q2 [1]),
    .C(\v0/z3/z4/z6/_01_ ),
    .X(\v0/z3/z4/z6/_03_ ));
 sky130_fd_sc_hd__lpflow_inputiso1p_1 \v0/z3/z4/z6/_25_  (.A(\v0/z3/z4/q3 [0]),
    .SLEEP(\v0/z3/z4/q2 [2]),
    .X(\v0/z3/z4/z6/_04_ ));
 sky130_fd_sc_hd__and2_0 \v0/z3/z4/z6/_26_  (.A(\v0/z3/z4/q3 [0]),
    .B(\v0/z3/z4/q2 [2]),
    .X(\v0/z3/z4/z6/_05_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z3/z4/z6/_27_  (.A(\v0/z3/z4/q3 [0]),
    .B(\v0/z3/z4/q2 [2]),
    .Y(\v0/z3/z4/z6/_06_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z3/z4/z6/_28_  (.A(\v0/z3/z4/z6/_04_ ),
    .B(\v0/z3/z4/z6/_06_ ),
    .Y(\v0/z3/z4/z6/_07_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z3/z4/z6/_29_  (.A(\v0/z3/z4/z6/_03_ ),
    .B(\v0/z3/z4/z6/_07_ ),
    .Y(\v0/z3/z4/q5 [2]));
 sky130_fd_sc_hd__nand2_1 \v0/z3/z4/z6/_30_  (.A(\v0/z3/z4/q3 [1]),
    .B(\v0/z3/z4/q2 [3]),
    .Y(\v0/z3/z4/z6/_08_ ));
 sky130_fd_sc_hd__xor2_1 \v0/z3/z4/z6/_31_  (.A(\v0/z3/z4/q3 [1]),
    .B(\v0/z3/z4/q2 [3]),
    .X(\v0/z3/z4/z6/_09_ ));
 sky130_fd_sc_hd__o21ai_0 \v0/z3/z4/z6/_32_  (.A1(\v0/z3/z4/z6/_03_ ),
    .A2(\v0/z3/z4/z6/_05_ ),
    .B1(\v0/z3/z4/z6/_04_ ),
    .Y(\v0/z3/z4/z6/_10_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z3/z4/z6/_33_  (.A(\v0/z3/z4/z6/_09_ ),
    .B(\v0/z3/z4/z6/_10_ ),
    .Y(\v0/z3/z4/q5 [3]));
 sky130_fd_sc_hd__nor2_1 \v0/z3/z4/z6/_34_  (.A(\v0/z3/z4/q3 [2]),
    .B(\v0/z3/z4/_03_ ),
    .Y(\v0/z3/z4/z6/_11_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z3/z4/z6/_35_  (.A(\v0/z3/z4/q3 [2]),
    .B(\v0/z3/z4/_03_ ),
    .Y(\v0/z3/z4/z6/_12_ ));
 sky130_fd_sc_hd__nand2b_1 \v0/z3/z4/z6/_36_  (.A_N(\v0/z3/z4/z6/_11_ ),
    .B(\v0/z3/z4/z6/_12_ ),
    .Y(\v0/z3/z4/z6/_13_ ));
 sky130_fd_sc_hd__o221ai_1 \v0/z3/z4/z6/_37_  (.A1(\v0/z3/z4/q3 [1]),
    .A2(\v0/z3/z4/q2 [3]),
    .B1(\v0/z3/z4/z6/_03_ ),
    .B2(\v0/z3/z4/z6/_05_ ),
    .C1(\v0/z3/z4/z6/_04_ ),
    .Y(\v0/z3/z4/z6/_14_ ));
 sky130_fd_sc_hd__a21oi_1 \v0/z3/z4/z6/_38_  (.A1(\v0/z3/z4/z6/_08_ ),
    .A2(\v0/z3/z4/z6/_14_ ),
    .B1(\v0/z3/z4/z6/_13_ ),
    .Y(\v0/z3/z4/z6/_15_ ));
 sky130_fd_sc_hd__and3_1 \v0/z3/z4/z6/_39_  (.A(\v0/z3/z4/z6/_08_ ),
    .B(\v0/z3/z4/z6/_13_ ),
    .C(\v0/z3/z4/z6/_14_ ),
    .X(\v0/z3/z4/z6/_16_ ));
 sky130_fd_sc_hd__nor2_1 \v0/z3/z4/z6/_40_  (.A(\v0/z3/z4/z6/_15_ ),
    .B(\v0/z3/z4/z6/_16_ ),
    .Y(\v0/z3/z4/q5 [4]));
 sky130_fd_sc_hd__xnor2_1 \v0/z3/z4/z6/_41_  (.A(\v0/z3/z4/q3 [3]),
    .B(\v0/z3/z4/_04_ ),
    .Y(\v0/z3/z4/z6/_17_ ));
 sky130_fd_sc_hd__a31oi_1 \v0/z3/z4/z6/_42_  (.A1(\v0/z3/z4/z6/_08_ ),
    .A2(\v0/z3/z4/z6/_12_ ),
    .A3(\v0/z3/z4/z6/_14_ ),
    .B1(\v0/z3/z4/z6/_11_ ),
    .Y(\v0/z3/z4/z6/_18_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z3/z4/z6/_43_  (.A(\v0/z3/z4/z6/_17_ ),
    .B(\v0/z3/z4/z6/_18_ ),
    .Y(\v0/z3/z4/q5 [5]));
 sky130_fd_sc_hd__maj3_1 \v0/z3/z4/z6/_44_  (.A(\v0/z3/z4/q3 [3]),
    .B(\v0/z3/z4/_04_ ),
    .C(\v0/z3/z4/z6/_18_ ),
    .X(\v0/z3/z4/z6/Cout ));
 sky130_fd_sc_hd__xnor2_1 \v0/z3/z4/z7/_19_  (.A(\v0/z3/z4/q5 [0]),
    .B(\v0/z3/z4/q4 [0]),
    .Y(\v0/z3/z4/z7/_00_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z3/z4/z7/_20_  (.A(\v0/z3/z4/_10_ ),
    .B(\v0/z3/z4/z7/_00_ ),
    .Y(\v0/z3/q3 [2]));
 sky130_fd_sc_hd__maj3_1 \v0/z3/z4/z7/_21_  (.A(\v0/z3/z4/q5 [0]),
    .B(\v0/z3/z4/q4 [0]),
    .C(\v0/z3/z4/_10_ ),
    .X(\v0/z3/z4/z7/_01_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z3/z4/z7/_22_  (.A(\v0/z3/z4/q5 [1]),
    .B(\v0/z3/z4/q4 [1]),
    .Y(\v0/z3/z4/z7/_02_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z3/z4/z7/_23_  (.A(\v0/z3/z4/z7/_01_ ),
    .B(\v0/z3/z4/z7/_02_ ),
    .Y(\v0/z3/q3 [3]));
 sky130_fd_sc_hd__maj3_1 \v0/z3/z4/z7/_24_  (.A(\v0/z3/z4/q5 [1]),
    .B(\v0/z3/z4/q4 [1]),
    .C(\v0/z3/z4/z7/_01_ ),
    .X(\v0/z3/z4/z7/_03_ ));
 sky130_fd_sc_hd__lpflow_inputiso1p_1 \v0/z3/z4/z7/_25_  (.A(\v0/z3/z4/q5 [2]),
    .SLEEP(\v0/z3/z4/q4 [2]),
    .X(\v0/z3/z4/z7/_04_ ));
 sky130_fd_sc_hd__and2_0 \v0/z3/z4/z7/_26_  (.A(\v0/z3/z4/q5 [2]),
    .B(\v0/z3/z4/q4 [2]),
    .X(\v0/z3/z4/z7/_05_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z3/z4/z7/_27_  (.A(\v0/z3/z4/q5 [2]),
    .B(\v0/z3/z4/q4 [2]),
    .Y(\v0/z3/z4/z7/_06_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z3/z4/z7/_28_  (.A(\v0/z3/z4/z7/_04_ ),
    .B(\v0/z3/z4/z7/_06_ ),
    .Y(\v0/z3/z4/z7/_07_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z3/z4/z7/_29_  (.A(\v0/z3/z4/z7/_03_ ),
    .B(\v0/z3/z4/z7/_07_ ),
    .Y(\v0/z3/q3 [4]));
 sky130_fd_sc_hd__nand2_1 \v0/z3/z4/z7/_30_  (.A(\v0/z3/z4/q5 [3]),
    .B(\v0/z3/z4/q4 [3]),
    .Y(\v0/z3/z4/z7/_08_ ));
 sky130_fd_sc_hd__xor2_1 \v0/z3/z4/z7/_31_  (.A(\v0/z3/z4/q5 [3]),
    .B(\v0/z3/z4/q4 [3]),
    .X(\v0/z3/z4/z7/_09_ ));
 sky130_fd_sc_hd__o21ai_0 \v0/z3/z4/z7/_32_  (.A1(\v0/z3/z4/z7/_03_ ),
    .A2(\v0/z3/z4/z7/_05_ ),
    .B1(\v0/z3/z4/z7/_04_ ),
    .Y(\v0/z3/z4/z7/_10_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z3/z4/z7/_33_  (.A(\v0/z3/z4/z7/_09_ ),
    .B(\v0/z3/z4/z7/_10_ ),
    .Y(\v0/z3/q3 [5]));
 sky130_fd_sc_hd__nor2_1 \v0/z3/z4/z7/_34_  (.A(\v0/z3/z4/q5 [4]),
    .B(\v0/z3/z4/_08_ ),
    .Y(\v0/z3/z4/z7/_11_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z3/z4/z7/_35_  (.A(\v0/z3/z4/q5 [4]),
    .B(\v0/z3/z4/_08_ ),
    .Y(\v0/z3/z4/z7/_12_ ));
 sky130_fd_sc_hd__nand2b_1 \v0/z3/z4/z7/_36_  (.A_N(\v0/z3/z4/z7/_11_ ),
    .B(\v0/z3/z4/z7/_12_ ),
    .Y(\v0/z3/z4/z7/_13_ ));
 sky130_fd_sc_hd__o221ai_1 \v0/z3/z4/z7/_37_  (.A1(\v0/z3/z4/q5 [3]),
    .A2(\v0/z3/z4/q4 [3]),
    .B1(\v0/z3/z4/z7/_03_ ),
    .B2(\v0/z3/z4/z7/_05_ ),
    .C1(\v0/z3/z4/z7/_04_ ),
    .Y(\v0/z3/z4/z7/_14_ ));
 sky130_fd_sc_hd__a21oi_1 \v0/z3/z4/z7/_38_  (.A1(\v0/z3/z4/z7/_08_ ),
    .A2(\v0/z3/z4/z7/_14_ ),
    .B1(\v0/z3/z4/z7/_13_ ),
    .Y(\v0/z3/z4/z7/_15_ ));
 sky130_fd_sc_hd__and3_1 \v0/z3/z4/z7/_39_  (.A(\v0/z3/z4/z7/_08_ ),
    .B(\v0/z3/z4/z7/_13_ ),
    .C(\v0/z3/z4/z7/_14_ ),
    .X(\v0/z3/z4/z7/_16_ ));
 sky130_fd_sc_hd__nor2_1 \v0/z3/z4/z7/_40_  (.A(\v0/z3/z4/z7/_15_ ),
    .B(\v0/z3/z4/z7/_16_ ),
    .Y(\v0/z3/q3 [6]));
 sky130_fd_sc_hd__xnor2_1 \v0/z3/z4/z7/_41_  (.A(\v0/z3/z4/q5 [5]),
    .B(\v0/z3/z4/_09_ ),
    .Y(\v0/z3/z4/z7/_17_ ));
 sky130_fd_sc_hd__a31oi_1 \v0/z3/z4/z7/_42_  (.A1(\v0/z3/z4/z7/_08_ ),
    .A2(\v0/z3/z4/z7/_12_ ),
    .A3(\v0/z3/z4/z7/_14_ ),
    .B1(\v0/z3/z4/z7/_11_ ),
    .Y(\v0/z3/z4/z7/_18_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z3/z4/z7/_43_  (.A(\v0/z3/z4/z7/_17_ ),
    .B(\v0/z3/z4/z7/_18_ ),
    .Y(\v0/z3/q3 [7]));
 sky130_fd_sc_hd__maj3_1 \v0/z3/z4/z7/_44_  (.A(\v0/z3/z4/q5 [5]),
    .B(\v0/z3/z4/_09_ ),
    .C(\v0/z3/z4/z7/_18_ ),
    .X(\v0/z3/z4/z7/Cout ));
 sky130_fd_sc_hd__xnor2_1 \v0/z3/z5/_27_  (.A(\v0/z3/q0 [4]),
    .B(\v0/z3/q1 [0]),
    .Y(\v0/z3/z5/_00_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z3/z5/_28_  (.A(\v0/z3/_04_ ),
    .B(\v0/z3/z5/_00_ ),
    .Y(\v0/z3/q4 [0]));
 sky130_fd_sc_hd__maj3_1 \v0/z3/z5/_29_  (.A(\v0/z3/q0 [4]),
    .B(\v0/z3/q1 [0]),
    .C(\v0/z3/_04_ ),
    .X(\v0/z3/z5/_01_ ));
 sky130_fd_sc_hd__lpflow_inputiso1p_1 \v0/z3/z5/_30_  (.A(\v0/z3/q0 [5]),
    .SLEEP(\v0/z3/q1 [1]),
    .X(\v0/z3/z5/_02_ ));
 sky130_fd_sc_hd__and2_0 \v0/z3/z5/_31_  (.A(\v0/z3/q0 [5]),
    .B(\v0/z3/q1 [1]),
    .X(\v0/z3/z5/_03_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z3/z5/_32_  (.A(\v0/z3/q0 [5]),
    .B(\v0/z3/q1 [1]),
    .Y(\v0/z3/z5/_04_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z3/z5/_33_  (.A(\v0/z3/z5/_02_ ),
    .B(\v0/z3/z5/_04_ ),
    .Y(\v0/z3/z5/_05_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z3/z5/_34_  (.A(\v0/z3/z5/_01_ ),
    .B(\v0/z3/z5/_05_ ),
    .Y(\v0/z3/q4 [1]));
 sky130_fd_sc_hd__nand2_1 \v0/z3/z5/_35_  (.A(\v0/z3/q0 [6]),
    .B(\v0/z3/q1 [2]),
    .Y(\v0/z3/z5/_06_ ));
 sky130_fd_sc_hd__xor2_1 \v0/z3/z5/_36_  (.A(\v0/z3/q0 [6]),
    .B(\v0/z3/q1 [2]),
    .X(\v0/z3/z5/_07_ ));
 sky130_fd_sc_hd__o21ai_0 \v0/z3/z5/_37_  (.A1(\v0/z3/z5/_01_ ),
    .A2(\v0/z3/z5/_03_ ),
    .B1(\v0/z3/z5/_02_ ),
    .Y(\v0/z3/z5/_08_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z3/z5/_38_  (.A(\v0/z3/z5/_07_ ),
    .B(\v0/z3/z5/_08_ ),
    .Y(\v0/z3/q4 [2]));
 sky130_fd_sc_hd__nor2_1 \v0/z3/z5/_39_  (.A(\v0/z3/q0 [7]),
    .B(\v0/z3/q1 [3]),
    .Y(\v0/z3/z5/_09_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z3/z5/_40_  (.A(\v0/z3/q0 [7]),
    .B(\v0/z3/q1 [3]),
    .Y(\v0/z3/z5/_10_ ));
 sky130_fd_sc_hd__nor2b_1 \v0/z3/z5/_41_  (.A(\v0/z3/z5/_09_ ),
    .B_N(\v0/z3/z5/_10_ ),
    .Y(\v0/z3/z5/_11_ ));
 sky130_fd_sc_hd__o221ai_1 \v0/z3/z5/_42_  (.A1(\v0/z3/q0 [6]),
    .A2(\v0/z3/q1 [2]),
    .B1(\v0/z3/z5/_01_ ),
    .B2(\v0/z3/z5/_03_ ),
    .C1(\v0/z3/z5/_02_ ),
    .Y(\v0/z3/z5/_12_ ));
 sky130_fd_sc_hd__and2_0 \v0/z3/z5/_43_  (.A(\v0/z3/z5/_06_ ),
    .B(\v0/z3/z5/_12_ ),
    .X(\v0/z3/z5/_13_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z3/z5/_44_  (.A(\v0/z3/z5/_11_ ),
    .B(\v0/z3/z5/_13_ ),
    .Y(\v0/z3/q4 [3]));
 sky130_fd_sc_hd__nor2_1 \v0/z3/z5/_45_  (.A(\v0/z3/_00_ ),
    .B(\v0/z3/q1 [4]),
    .Y(\v0/z3/z5/_14_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z3/z5/_46_  (.A(\v0/z3/_00_ ),
    .B(\v0/z3/q1 [4]),
    .Y(\v0/z3/z5/_15_ ));
 sky130_fd_sc_hd__nand2b_1 \v0/z3/z5/_47_  (.A_N(\v0/z3/z5/_14_ ),
    .B(\v0/z3/z5/_15_ ),
    .Y(\v0/z3/z5/_16_ ));
 sky130_fd_sc_hd__a21oi_1 \v0/z3/z5/_48_  (.A1(\v0/z3/z5/_10_ ),
    .A2(\v0/z3/z5/_13_ ),
    .B1(\v0/z3/z5/_09_ ),
    .Y(\v0/z3/z5/_17_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z3/z5/_49_  (.A(\v0/z3/z5/_16_ ),
    .B(\v0/z3/z5/_17_ ),
    .Y(\v0/z3/q4 [4]));
 sky130_fd_sc_hd__a311o_1 \v0/z3/z5/_50_  (.A1(\v0/z3/z5/_06_ ),
    .A2(\v0/z3/z5/_10_ ),
    .A3(\v0/z3/z5/_12_ ),
    .B1(\v0/z3/z5/_14_ ),
    .C1(\v0/z3/z5/_09_ ),
    .X(\v0/z3/z5/_18_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z3/z5/_51_  (.A(\v0/z3/z5/_15_ ),
    .B(\v0/z3/z5/_18_ ),
    .Y(\v0/z3/z5/_19_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z3/z5/_52_  (.A(\v0/z3/_01_ ),
    .B(\v0/z3/q1 [5]),
    .Y(\v0/z3/z5/_20_ ));
 sky130_fd_sc_hd__nor2_1 \v0/z3/z5/_53_  (.A(\v0/z3/_01_ ),
    .B(\v0/z3/q1 [5]),
    .Y(\v0/z3/z5/_21_ ));
 sky130_fd_sc_hd__a31oi_1 \v0/z3/z5/_54_  (.A1(\v0/z3/z5/_15_ ),
    .A2(\v0/z3/z5/_18_ ),
    .A3(\v0/z3/z5/_20_ ),
    .B1(\v0/z3/z5/_21_ ),
    .Y(\v0/z3/z5/_22_ ));
 sky130_fd_sc_hd__a21bo_1 \v0/z3/z5/_55_  (.A1(\v0/z3/z5/_20_ ),
    .A2(\v0/z3/z5/_22_ ),
    .B1_N(\v0/z3/z5/_19_ ),
    .X(\v0/z3/z5/_23_ ));
 sky130_fd_sc_hd__o21ai_0 \v0/z3/z5/_56_  (.A1(\v0/z3/z5/_21_ ),
    .A2(\v0/z3/z5/_22_ ),
    .B1(\v0/z3/z5/_23_ ),
    .Y(\v0/z3/q4 [5]));
 sky130_fd_sc_hd__xnor2_1 \v0/z3/z5/_57_  (.A(\v0/z3/_02_ ),
    .B(\v0/z3/q1 [6]),
    .Y(\v0/z3/z5/_24_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z3/z5/_58_  (.A(\v0/z3/z5/_22_ ),
    .B(\v0/z3/z5/_24_ ),
    .Y(\v0/z3/q4 [6]));
 sky130_fd_sc_hd__xnor2_1 \v0/z3/z5/_59_  (.A(\v0/z3/_03_ ),
    .B(\v0/z3/q1 [7]),
    .Y(\v0/z3/z5/_25_ ));
 sky130_fd_sc_hd__maj3_1 \v0/z3/z5/_60_  (.A(\v0/z3/_02_ ),
    .B(\v0/z3/q1 [6]),
    .C(\v0/z3/z5/_22_ ),
    .X(\v0/z3/z5/_26_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z3/z5/_61_  (.A(\v0/z3/z5/_25_ ),
    .B(\v0/z3/z5/_26_ ),
    .Y(\v0/z3/q4 [7]));
 sky130_fd_sc_hd__maj3_1 \v0/z3/z5/_62_  (.A(\v0/z3/_03_ ),
    .B(\v0/z3/q1 [7]),
    .C(\v0/z3/z5/_26_ ),
    .X(\v0/z3/z5/Cout ));
 sky130_fd_sc_hd__xnor2_1 \v0/z3/z6/_050_  (.A(\v0/z3/_09_ ),
    .B(\v0/z3/q2 [0]),
    .Y(\v0/z3/z6/_000_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z3/z6/_051_  (.A(\v0/z3/_13_ ),
    .B(\v0/z3/z6/_000_ ),
    .Y(\v0/z3/q5 [0]));
 sky130_fd_sc_hd__maj3_1 \v0/z3/z6/_052_  (.A(\v0/z3/_09_ ),
    .B(\v0/z3/q2 [0]),
    .C(\v0/z3/_13_ ),
    .X(\v0/z3/z6/_001_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z3/z6/_053_  (.A(\v0/z3/_10_ ),
    .B(\v0/z3/q2 [1]),
    .Y(\v0/z3/z6/_002_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z3/z6/_054_  (.A(\v0/z3/z6/_001_ ),
    .B(\v0/z3/z6/_002_ ),
    .Y(\v0/z3/q5 [1]));
 sky130_fd_sc_hd__maj3_1 \v0/z3/z6/_055_  (.A(\v0/z3/_10_ ),
    .B(\v0/z3/q2 [1]),
    .C(\v0/z3/z6/_001_ ),
    .X(\v0/z3/z6/_003_ ));
 sky130_fd_sc_hd__lpflow_inputiso1p_1 \v0/z3/z6/_056_  (.A(\v0/z3/_11_ ),
    .SLEEP(\v0/z3/q2 [2]),
    .X(\v0/z3/z6/_004_ ));
 sky130_fd_sc_hd__and2_0 \v0/z3/z6/_057_  (.A(\v0/z3/_11_ ),
    .B(\v0/z3/q2 [2]),
    .X(\v0/z3/z6/_005_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z3/z6/_058_  (.A(\v0/z3/_11_ ),
    .B(\v0/z3/q2 [2]),
    .Y(\v0/z3/z6/_006_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z3/z6/_059_  (.A(\v0/z3/z6/_004_ ),
    .B(\v0/z3/z6/_006_ ),
    .Y(\v0/z3/z6/_007_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z3/z6/_060_  (.A(\v0/z3/z6/_003_ ),
    .B(\v0/z3/z6/_007_ ),
    .Y(\v0/z3/q5 [2]));
 sky130_fd_sc_hd__nor2_1 \v0/z3/z6/_061_  (.A(\v0/z3/_12_ ),
    .B(\v0/z3/q2 [3]),
    .Y(\v0/z3/z6/_008_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z3/z6/_062_  (.A(\v0/z3/_12_ ),
    .B(\v0/z3/q2 [3]),
    .Y(\v0/z3/z6/_009_ ));
 sky130_fd_sc_hd__clkinv_1 \v0/z3/z6/_063_  (.A(\v0/z3/z6/_009_ ),
    .Y(\v0/z3/z6/_010_ ));
 sky130_fd_sc_hd__nor2_1 \v0/z3/z6/_064_  (.A(\v0/z3/z6/_008_ ),
    .B(\v0/z3/z6/_010_ ),
    .Y(\v0/z3/z6/_011_ ));
 sky130_fd_sc_hd__o21ai_0 \v0/z3/z6/_065_  (.A1(\v0/z3/z6/_003_ ),
    .A2(\v0/z3/z6/_005_ ),
    .B1(\v0/z3/z6/_004_ ),
    .Y(\v0/z3/z6/_012_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z3/z6/_066_  (.A(\v0/z3/z6/_011_ ),
    .B(\v0/z3/z6/_012_ ),
    .Y(\v0/z3/q5 [3]));
 sky130_fd_sc_hd__lpflow_inputiso1p_1 \v0/z3/z6/_067_  (.A(\v0/z3/q3 [0]),
    .SLEEP(\v0/z3/q2 [4]),
    .X(\v0/z3/z6/_013_ ));
 sky130_fd_sc_hd__and2_0 \v0/z3/z6/_068_  (.A(\v0/z3/q3 [0]),
    .B(\v0/z3/q2 [4]),
    .X(\v0/z3/z6/_014_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z3/z6/_069_  (.A(\v0/z3/q3 [0]),
    .B(\v0/z3/q2 [4]),
    .Y(\v0/z3/z6/_015_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z3/z6/_070_  (.A(\v0/z3/z6/_013_ ),
    .B(\v0/z3/z6/_015_ ),
    .Y(\v0/z3/z6/_016_ ));
 sky130_fd_sc_hd__o221a_1 \v0/z3/z6/_071_  (.A1(\v0/z3/_12_ ),
    .A2(\v0/z3/q2 [3]),
    .B1(\v0/z3/z6/_003_ ),
    .B2(\v0/z3/z6/_005_ ),
    .C1(\v0/z3/z6/_004_ ),
    .X(\v0/z3/z6/_017_ ));
 sky130_fd_sc_hd__a21oi_1 \v0/z3/z6/_072_  (.A1(\v0/z3/z6/_009_ ),
    .A2(\v0/z3/z6/_012_ ),
    .B1(\v0/z3/z6/_008_ ),
    .Y(\v0/z3/z6/_018_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z3/z6/_073_  (.A(\v0/z3/z6/_016_ ),
    .B(\v0/z3/z6/_018_ ),
    .Y(\v0/z3/q5 [4]));
 sky130_fd_sc_hd__lpflow_inputiso1p_1 \v0/z3/z6/_074_  (.A(\v0/z3/q3 [1]),
    .SLEEP(\v0/z3/q2 [5]),
    .X(\v0/z3/z6/_019_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z3/z6/_075_  (.A(\v0/z3/q3 [1]),
    .B(\v0/z3/q2 [5]),
    .Y(\v0/z3/z6/_020_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z3/z6/_076_  (.A(\v0/z3/z6/_019_ ),
    .B(\v0/z3/z6/_020_ ),
    .Y(\v0/z3/z6/_021_ ));
 sky130_fd_sc_hd__o21ai_0 \v0/z3/z6/_077_  (.A1(\v0/z3/z6/_014_ ),
    .A2(\v0/z3/z6/_018_ ),
    .B1(\v0/z3/z6/_013_ ),
    .Y(\v0/z3/z6/_022_ ));
 sky130_fd_sc_hd__xor2_1 \v0/z3/z6/_078_  (.A(\v0/z3/z6/_021_ ),
    .B(\v0/z3/z6/_022_ ),
    .X(\v0/z3/q5 [5]));
 sky130_fd_sc_hd__nor2_1 \v0/z3/z6/_079_  (.A(\v0/z3/q3 [2]),
    .B(\v0/z3/q2 [6]),
    .Y(\v0/z3/z6/_023_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z3/z6/_080_  (.A(\v0/z3/q3 [2]),
    .B(\v0/z3/q2 [6]),
    .Y(\v0/z3/z6/_024_ ));
 sky130_fd_sc_hd__nor2b_1 \v0/z3/z6/_081_  (.A(\v0/z3/z6/_023_ ),
    .B_N(\v0/z3/z6/_024_ ),
    .Y(\v0/z3/z6/_025_ ));
 sky130_fd_sc_hd__o311ai_0 \v0/z3/z6/_082_  (.A1(\v0/z3/z6/_010_ ),
    .A2(\v0/z3/z6/_014_ ),
    .A3(\v0/z3/z6/_017_ ),
    .B1(\v0/z3/z6/_019_ ),
    .C1(\v0/z3/z6/_013_ ),
    .Y(\v0/z3/z6/_026_ ));
 sky130_fd_sc_hd__and2_0 \v0/z3/z6/_083_  (.A(\v0/z3/z6/_020_ ),
    .B(\v0/z3/z6/_026_ ),
    .X(\v0/z3/z6/_027_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z3/z6/_084_  (.A(\v0/z3/z6/_025_ ),
    .B(\v0/z3/z6/_027_ ),
    .Y(\v0/z3/q5 [6]));
 sky130_fd_sc_hd__nor2_1 \v0/z3/z6/_085_  (.A(\v0/z3/q3 [3]),
    .B(\v0/z3/q2 [7]),
    .Y(\v0/z3/z6/_028_ ));
 sky130_fd_sc_hd__and2_0 \v0/z3/z6/_086_  (.A(\v0/z3/q3 [3]),
    .B(\v0/z3/q2 [7]),
    .X(\v0/z3/z6/_029_ ));
 sky130_fd_sc_hd__nor2_1 \v0/z3/z6/_087_  (.A(\v0/z3/z6/_028_ ),
    .B(\v0/z3/z6/_029_ ),
    .Y(\v0/z3/z6/_030_ ));
 sky130_fd_sc_hd__a21oi_1 \v0/z3/z6/_088_  (.A1(\v0/z3/z6/_024_ ),
    .A2(\v0/z3/z6/_027_ ),
    .B1(\v0/z3/z6/_023_ ),
    .Y(\v0/z3/z6/_031_ ));
 sky130_fd_sc_hd__xor2_1 \v0/z3/z6/_089_  (.A(\v0/z3/z6/_030_ ),
    .B(\v0/z3/z6/_031_ ),
    .X(\v0/z3/q5 [7]));
 sky130_fd_sc_hd__lpflow_inputiso1p_1 \v0/z3/z6/_090_  (.A(\v0/z3/q3 [4]),
    .SLEEP(\v0/z3/_05_ ),
    .X(\v0/z3/z6/_032_ ));
 sky130_fd_sc_hd__and2_0 \v0/z3/z6/_091_  (.A(\v0/z3/q3 [4]),
    .B(\v0/z3/_05_ ),
    .X(\v0/z3/z6/_033_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z3/z6/_092_  (.A(\v0/z3/q3 [4]),
    .B(\v0/z3/_05_ ),
    .Y(\v0/z3/z6/_034_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z3/z6/_093_  (.A(\v0/z3/z6/_032_ ),
    .B(\v0/z3/z6/_034_ ),
    .Y(\v0/z3/z6/_035_ ));
 sky130_fd_sc_hd__a311oi_1 \v0/z3/z6/_094_  (.A1(\v0/z3/z6/_020_ ),
    .A2(\v0/z3/z6/_024_ ),
    .A3(\v0/z3/z6/_026_ ),
    .B1(\v0/z3/z6/_028_ ),
    .C1(\v0/z3/z6/_023_ ),
    .Y(\v0/z3/z6/_036_ ));
 sky130_fd_sc_hd__lpflow_inputiso1p_1 \v0/z3/z6/_095_  (.A(\v0/z3/z6/_029_ ),
    .SLEEP(\v0/z3/z6/_036_ ),
    .X(\v0/z3/z6/_037_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z3/z6/_096_  (.A(\v0/z3/z6/_035_ ),
    .B(\v0/z3/z6/_037_ ),
    .Y(\v0/z3/q5 [8]));
 sky130_fd_sc_hd__lpflow_inputiso1p_1 \v0/z3/z6/_097_  (.A(\v0/z3/q3 [5]),
    .SLEEP(\v0/z3/_06_ ),
    .X(\v0/z3/z6/_038_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z3/z6/_098_  (.A(\v0/z3/q3 [5]),
    .B(\v0/z3/_06_ ),
    .Y(\v0/z3/z6/_039_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z3/z6/_099_  (.A(\v0/z3/z6/_038_ ),
    .B(\v0/z3/z6/_039_ ),
    .Y(\v0/z3/z6/_040_ ));
 sky130_fd_sc_hd__o21ai_0 \v0/z3/z6/_100_  (.A1(\v0/z3/z6/_033_ ),
    .A2(\v0/z3/z6/_037_ ),
    .B1(\v0/z3/z6/_032_ ),
    .Y(\v0/z3/z6/_041_ ));
 sky130_fd_sc_hd__xor2_1 \v0/z3/z6/_101_  (.A(\v0/z3/z6/_040_ ),
    .B(\v0/z3/z6/_041_ ),
    .X(\v0/z3/q5 [9]));
 sky130_fd_sc_hd__nor2_1 \v0/z3/z6/_102_  (.A(\v0/z3/q3 [6]),
    .B(\v0/z3/_07_ ),
    .Y(\v0/z3/z6/_042_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z3/z6/_103_  (.A(\v0/z3/q3 [6]),
    .B(\v0/z3/_07_ ),
    .Y(\v0/z3/z6/_043_ ));
 sky130_fd_sc_hd__nand2b_1 \v0/z3/z6/_104_  (.A_N(\v0/z3/z6/_042_ ),
    .B(\v0/z3/z6/_043_ ),
    .Y(\v0/z3/z6/_044_ ));
 sky130_fd_sc_hd__o311ai_0 \v0/z3/z6/_105_  (.A1(\v0/z3/z6/_029_ ),
    .A2(\v0/z3/z6/_033_ ),
    .A3(\v0/z3/z6/_036_ ),
    .B1(\v0/z3/z6/_038_ ),
    .C1(\v0/z3/z6/_032_ ),
    .Y(\v0/z3/z6/_045_ ));
 sky130_fd_sc_hd__a21oi_1 \v0/z3/z6/_106_  (.A1(\v0/z3/z6/_039_ ),
    .A2(\v0/z3/z6/_045_ ),
    .B1(\v0/z3/z6/_044_ ),
    .Y(\v0/z3/z6/_046_ ));
 sky130_fd_sc_hd__and3_1 \v0/z3/z6/_107_  (.A(\v0/z3/z6/_039_ ),
    .B(\v0/z3/z6/_044_ ),
    .C(\v0/z3/z6/_045_ ),
    .X(\v0/z3/z6/_047_ ));
 sky130_fd_sc_hd__nor2_1 \v0/z3/z6/_108_  (.A(\v0/z3/z6/_046_ ),
    .B(\v0/z3/z6/_047_ ),
    .Y(\v0/z3/q5 [10]));
 sky130_fd_sc_hd__xnor2_1 \v0/z3/z6/_109_  (.A(\v0/z3/q3 [7]),
    .B(\v0/z3/_08_ ),
    .Y(\v0/z3/z6/_048_ ));
 sky130_fd_sc_hd__a31oi_1 \v0/z3/z6/_110_  (.A1(\v0/z3/z6/_039_ ),
    .A2(\v0/z3/z6/_043_ ),
    .A3(\v0/z3/z6/_045_ ),
    .B1(\v0/z3/z6/_042_ ),
    .Y(\v0/z3/z6/_049_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z3/z6/_111_  (.A(\v0/z3/z6/_048_ ),
    .B(\v0/z3/z6/_049_ ),
    .Y(\v0/z3/q5 [11]));
 sky130_fd_sc_hd__maj3_1 \v0/z3/z6/_112_  (.A(\v0/z3/q3 [7]),
    .B(\v0/z3/_08_ ),
    .C(\v0/z3/z6/_049_ ),
    .X(\v0/z3/z6/Cout ));
 sky130_fd_sc_hd__xnor2_1 \v0/z3/z7/_050_  (.A(\v0/z3/q5 [0]),
    .B(\v0/z3/q4 [0]),
    .Y(\v0/z3/z7/_000_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z3/z7/_051_  (.A(\v0/z3/_18_ ),
    .B(\v0/z3/z7/_000_ ),
    .Y(\v0/q2 [4]));
 sky130_fd_sc_hd__maj3_1 \v0/z3/z7/_052_  (.A(\v0/z3/q5 [0]),
    .B(\v0/z3/q4 [0]),
    .C(\v0/z3/_18_ ),
    .X(\v0/z3/z7/_001_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z3/z7/_053_  (.A(\v0/z3/q5 [1]),
    .B(\v0/z3/q4 [1]),
    .Y(\v0/z3/z7/_002_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z3/z7/_054_  (.A(\v0/z3/z7/_001_ ),
    .B(\v0/z3/z7/_002_ ),
    .Y(\v0/q2 [5]));
 sky130_fd_sc_hd__maj3_1 \v0/z3/z7/_055_  (.A(\v0/z3/q5 [1]),
    .B(\v0/z3/q4 [1]),
    .C(\v0/z3/z7/_001_ ),
    .X(\v0/z3/z7/_003_ ));
 sky130_fd_sc_hd__lpflow_inputiso1p_1 \v0/z3/z7/_056_  (.A(\v0/z3/q5 [2]),
    .SLEEP(\v0/z3/q4 [2]),
    .X(\v0/z3/z7/_004_ ));
 sky130_fd_sc_hd__and2_0 \v0/z3/z7/_057_  (.A(\v0/z3/q5 [2]),
    .B(\v0/z3/q4 [2]),
    .X(\v0/z3/z7/_005_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z3/z7/_058_  (.A(\v0/z3/q5 [2]),
    .B(\v0/z3/q4 [2]),
    .Y(\v0/z3/z7/_006_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z3/z7/_059_  (.A(\v0/z3/z7/_004_ ),
    .B(\v0/z3/z7/_006_ ),
    .Y(\v0/z3/z7/_007_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z3/z7/_060_  (.A(\v0/z3/z7/_003_ ),
    .B(\v0/z3/z7/_007_ ),
    .Y(\v0/q2 [6]));
 sky130_fd_sc_hd__nor2_1 \v0/z3/z7/_061_  (.A(\v0/z3/q5 [3]),
    .B(\v0/z3/q4 [3]),
    .Y(\v0/z3/z7/_008_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z3/z7/_062_  (.A(\v0/z3/q5 [3]),
    .B(\v0/z3/q4 [3]),
    .Y(\v0/z3/z7/_009_ ));
 sky130_fd_sc_hd__clkinv_1 \v0/z3/z7/_063_  (.A(\v0/z3/z7/_009_ ),
    .Y(\v0/z3/z7/_010_ ));
 sky130_fd_sc_hd__nor2_1 \v0/z3/z7/_064_  (.A(\v0/z3/z7/_008_ ),
    .B(\v0/z3/z7/_010_ ),
    .Y(\v0/z3/z7/_011_ ));
 sky130_fd_sc_hd__o21ai_0 \v0/z3/z7/_065_  (.A1(\v0/z3/z7/_003_ ),
    .A2(\v0/z3/z7/_005_ ),
    .B1(\v0/z3/z7/_004_ ),
    .Y(\v0/z3/z7/_012_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z3/z7/_066_  (.A(\v0/z3/z7/_011_ ),
    .B(\v0/z3/z7/_012_ ),
    .Y(\v0/q2 [7]));
 sky130_fd_sc_hd__lpflow_inputiso1p_1 \v0/z3/z7/_067_  (.A(\v0/z3/q5 [4]),
    .SLEEP(\v0/z3/q4 [4]),
    .X(\v0/z3/z7/_013_ ));
 sky130_fd_sc_hd__and2_0 \v0/z3/z7/_068_  (.A(\v0/z3/q5 [4]),
    .B(\v0/z3/q4 [4]),
    .X(\v0/z3/z7/_014_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z3/z7/_069_  (.A(\v0/z3/q5 [4]),
    .B(\v0/z3/q4 [4]),
    .Y(\v0/z3/z7/_015_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z3/z7/_070_  (.A(\v0/z3/z7/_013_ ),
    .B(\v0/z3/z7/_015_ ),
    .Y(\v0/z3/z7/_016_ ));
 sky130_fd_sc_hd__o221a_1 \v0/z3/z7/_071_  (.A1(\v0/z3/q5 [3]),
    .A2(\v0/z3/q4 [3]),
    .B1(\v0/z3/z7/_003_ ),
    .B2(\v0/z3/z7/_005_ ),
    .C1(\v0/z3/z7/_004_ ),
    .X(\v0/z3/z7/_017_ ));
 sky130_fd_sc_hd__a21oi_1 \v0/z3/z7/_072_  (.A1(\v0/z3/z7/_009_ ),
    .A2(\v0/z3/z7/_012_ ),
    .B1(\v0/z3/z7/_008_ ),
    .Y(\v0/z3/z7/_018_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z3/z7/_073_  (.A(\v0/z3/z7/_016_ ),
    .B(\v0/z3/z7/_018_ ),
    .Y(\v0/q2 [8]));
 sky130_fd_sc_hd__lpflow_inputiso1p_1 \v0/z3/z7/_074_  (.A(\v0/z3/q5 [5]),
    .SLEEP(\v0/z3/q4 [5]),
    .X(\v0/z3/z7/_019_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z3/z7/_075_  (.A(\v0/z3/q5 [5]),
    .B(\v0/z3/q4 [5]),
    .Y(\v0/z3/z7/_020_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z3/z7/_076_  (.A(\v0/z3/z7/_019_ ),
    .B(\v0/z3/z7/_020_ ),
    .Y(\v0/z3/z7/_021_ ));
 sky130_fd_sc_hd__o21ai_0 \v0/z3/z7/_077_  (.A1(\v0/z3/z7/_014_ ),
    .A2(\v0/z3/z7/_018_ ),
    .B1(\v0/z3/z7/_013_ ),
    .Y(\v0/z3/z7/_022_ ));
 sky130_fd_sc_hd__xor2_1 \v0/z3/z7/_078_  (.A(\v0/z3/z7/_021_ ),
    .B(\v0/z3/z7/_022_ ),
    .X(\v0/q2 [9]));
 sky130_fd_sc_hd__nor2_1 \v0/z3/z7/_079_  (.A(\v0/z3/q5 [6]),
    .B(\v0/z3/q4 [6]),
    .Y(\v0/z3/z7/_023_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z3/z7/_080_  (.A(\v0/z3/q5 [6]),
    .B(\v0/z3/q4 [6]),
    .Y(\v0/z3/z7/_024_ ));
 sky130_fd_sc_hd__nor2b_1 \v0/z3/z7/_081_  (.A(\v0/z3/z7/_023_ ),
    .B_N(\v0/z3/z7/_024_ ),
    .Y(\v0/z3/z7/_025_ ));
 sky130_fd_sc_hd__o311ai_0 \v0/z3/z7/_082_  (.A1(\v0/z3/z7/_010_ ),
    .A2(\v0/z3/z7/_014_ ),
    .A3(\v0/z3/z7/_017_ ),
    .B1(\v0/z3/z7/_019_ ),
    .C1(\v0/z3/z7/_013_ ),
    .Y(\v0/z3/z7/_026_ ));
 sky130_fd_sc_hd__and2_0 \v0/z3/z7/_083_  (.A(\v0/z3/z7/_020_ ),
    .B(\v0/z3/z7/_026_ ),
    .X(\v0/z3/z7/_027_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z3/z7/_084_  (.A(\v0/z3/z7/_025_ ),
    .B(\v0/z3/z7/_027_ ),
    .Y(\v0/q2 [10]));
 sky130_fd_sc_hd__nor2_1 \v0/z3/z7/_085_  (.A(\v0/z3/q5 [7]),
    .B(\v0/z3/q4 [7]),
    .Y(\v0/z3/z7/_028_ ));
 sky130_fd_sc_hd__and2_0 \v0/z3/z7/_086_  (.A(\v0/z3/q5 [7]),
    .B(\v0/z3/q4 [7]),
    .X(\v0/z3/z7/_029_ ));
 sky130_fd_sc_hd__nor2_1 \v0/z3/z7/_087_  (.A(\v0/z3/z7/_028_ ),
    .B(\v0/z3/z7/_029_ ),
    .Y(\v0/z3/z7/_030_ ));
 sky130_fd_sc_hd__a21oi_1 \v0/z3/z7/_088_  (.A1(\v0/z3/z7/_024_ ),
    .A2(\v0/z3/z7/_027_ ),
    .B1(\v0/z3/z7/_023_ ),
    .Y(\v0/z3/z7/_031_ ));
 sky130_fd_sc_hd__xor2_1 \v0/z3/z7/_089_  (.A(\v0/z3/z7/_030_ ),
    .B(\v0/z3/z7/_031_ ),
    .X(\v0/q2 [11]));
 sky130_fd_sc_hd__lpflow_inputiso1p_1 \v0/z3/z7/_090_  (.A(\v0/z3/q5 [8]),
    .SLEEP(\v0/z3/_14_ ),
    .X(\v0/z3/z7/_032_ ));
 sky130_fd_sc_hd__and2_0 \v0/z3/z7/_091_  (.A(\v0/z3/q5 [8]),
    .B(\v0/z3/_14_ ),
    .X(\v0/z3/z7/_033_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z3/z7/_092_  (.A(\v0/z3/q5 [8]),
    .B(\v0/z3/_14_ ),
    .Y(\v0/z3/z7/_034_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z3/z7/_093_  (.A(\v0/z3/z7/_032_ ),
    .B(\v0/z3/z7/_034_ ),
    .Y(\v0/z3/z7/_035_ ));
 sky130_fd_sc_hd__a311oi_1 \v0/z3/z7/_094_  (.A1(\v0/z3/z7/_020_ ),
    .A2(\v0/z3/z7/_024_ ),
    .A3(\v0/z3/z7/_026_ ),
    .B1(\v0/z3/z7/_028_ ),
    .C1(\v0/z3/z7/_023_ ),
    .Y(\v0/z3/z7/_036_ ));
 sky130_fd_sc_hd__lpflow_inputiso1p_1 \v0/z3/z7/_095_  (.A(\v0/z3/z7/_029_ ),
    .SLEEP(\v0/z3/z7/_036_ ),
    .X(\v0/z3/z7/_037_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z3/z7/_096_  (.A(\v0/z3/z7/_035_ ),
    .B(\v0/z3/z7/_037_ ),
    .Y(\v0/q2 [12]));
 sky130_fd_sc_hd__lpflow_inputiso1p_1 \v0/z3/z7/_097_  (.A(\v0/z3/q5 [9]),
    .SLEEP(\v0/z3/_15_ ),
    .X(\v0/z3/z7/_038_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z3/z7/_098_  (.A(\v0/z3/q5 [9]),
    .B(\v0/z3/_15_ ),
    .Y(\v0/z3/z7/_039_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z3/z7/_099_  (.A(\v0/z3/z7/_038_ ),
    .B(\v0/z3/z7/_039_ ),
    .Y(\v0/z3/z7/_040_ ));
 sky130_fd_sc_hd__o21ai_0 \v0/z3/z7/_100_  (.A1(\v0/z3/z7/_033_ ),
    .A2(\v0/z3/z7/_037_ ),
    .B1(\v0/z3/z7/_032_ ),
    .Y(\v0/z3/z7/_041_ ));
 sky130_fd_sc_hd__xor2_1 \v0/z3/z7/_101_  (.A(\v0/z3/z7/_040_ ),
    .B(\v0/z3/z7/_041_ ),
    .X(\v0/q2 [13]));
 sky130_fd_sc_hd__nor2_1 \v0/z3/z7/_102_  (.A(\v0/z3/q5 [10]),
    .B(\v0/z3/_16_ ),
    .Y(\v0/z3/z7/_042_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z3/z7/_103_  (.A(\v0/z3/q5 [10]),
    .B(\v0/z3/_16_ ),
    .Y(\v0/z3/z7/_043_ ));
 sky130_fd_sc_hd__nand2b_1 \v0/z3/z7/_104_  (.A_N(\v0/z3/z7/_042_ ),
    .B(\v0/z3/z7/_043_ ),
    .Y(\v0/z3/z7/_044_ ));
 sky130_fd_sc_hd__o311ai_0 \v0/z3/z7/_105_  (.A1(\v0/z3/z7/_029_ ),
    .A2(\v0/z3/z7/_033_ ),
    .A3(\v0/z3/z7/_036_ ),
    .B1(\v0/z3/z7/_038_ ),
    .C1(\v0/z3/z7/_032_ ),
    .Y(\v0/z3/z7/_045_ ));
 sky130_fd_sc_hd__a21oi_1 \v0/z3/z7/_106_  (.A1(\v0/z3/z7/_039_ ),
    .A2(\v0/z3/z7/_045_ ),
    .B1(\v0/z3/z7/_044_ ),
    .Y(\v0/z3/z7/_046_ ));
 sky130_fd_sc_hd__and3_1 \v0/z3/z7/_107_  (.A(\v0/z3/z7/_039_ ),
    .B(\v0/z3/z7/_044_ ),
    .C(\v0/z3/z7/_045_ ),
    .X(\v0/z3/z7/_047_ ));
 sky130_fd_sc_hd__nor2_1 \v0/z3/z7/_108_  (.A(\v0/z3/z7/_046_ ),
    .B(\v0/z3/z7/_047_ ),
    .Y(\v0/q2 [14]));
 sky130_fd_sc_hd__xnor2_1 \v0/z3/z7/_109_  (.A(\v0/z3/q5 [11]),
    .B(\v0/z3/_17_ ),
    .Y(\v0/z3/z7/_048_ ));
 sky130_fd_sc_hd__a31oi_1 \v0/z3/z7/_110_  (.A1(\v0/z3/z7/_039_ ),
    .A2(\v0/z3/z7/_043_ ),
    .A3(\v0/z3/z7/_045_ ),
    .B1(\v0/z3/z7/_042_ ),
    .Y(\v0/z3/z7/_049_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z3/z7/_111_  (.A(\v0/z3/z7/_048_ ),
    .B(\v0/z3/z7/_049_ ),
    .Y(\v0/q2 [15]));
 sky130_fd_sc_hd__maj3_1 \v0/z3/z7/_112_  (.A(\v0/z3/q5 [11]),
    .B(\v0/z3/_17_ ),
    .C(\v0/z3/z7/_049_ ),
    .X(\v0/z3/z7/Cout ));
 sky130_fd_sc_hd__conb_1 \v0/z4/_19_  (.LO(\v0/z4/_00_ ));
 sky130_fd_sc_hd__conb_1 \v0/z4/_20_  (.LO(\v0/z4/_01_ ));
 sky130_fd_sc_hd__conb_1 \v0/z4/_21_  (.LO(\v0/z4/_02_ ));
 sky130_fd_sc_hd__conb_1 \v0/z4/_22_  (.LO(\v0/z4/_03_ ));
 sky130_fd_sc_hd__conb_1 \v0/z4/_23_  (.LO(\v0/z4/_04_ ));
 sky130_fd_sc_hd__conb_1 \v0/z4/_24_  (.LO(\v0/z4/_05_ ));
 sky130_fd_sc_hd__conb_1 \v0/z4/_25_  (.LO(\v0/z4/_06_ ));
 sky130_fd_sc_hd__conb_1 \v0/z4/_26_  (.LO(\v0/z4/_07_ ));
 sky130_fd_sc_hd__conb_1 \v0/z4/_27_  (.LO(\v0/z4/_08_ ));
 sky130_fd_sc_hd__conb_1 \v0/z4/_28_  (.LO(\v0/z4/_09_ ));
 sky130_fd_sc_hd__conb_1 \v0/z4/_29_  (.LO(\v0/z4/_10_ ));
 sky130_fd_sc_hd__conb_1 \v0/z4/_30_  (.LO(\v0/z4/_11_ ));
 sky130_fd_sc_hd__conb_1 \v0/z4/_31_  (.LO(\v0/z4/_12_ ));
 sky130_fd_sc_hd__conb_1 \v0/z4/_32_  (.LO(\v0/z4/_13_ ));
 sky130_fd_sc_hd__conb_1 \v0/z4/_33_  (.LO(\v0/z4/_14_ ));
 sky130_fd_sc_hd__conb_1 \v0/z4/_34_  (.LO(\v0/z4/_15_ ));
 sky130_fd_sc_hd__conb_1 \v0/z4/_35_  (.LO(\v0/z4/_16_ ));
 sky130_fd_sc_hd__conb_1 \v0/z4/_36_  (.LO(\v0/z4/_17_ ));
 sky130_fd_sc_hd__conb_1 \v0/z4/_37_  (.LO(\v0/z4/_18_ ));
 sky130_fd_sc_hd__conb_1 \v0/z4/z1/_11_  (.LO(\v0/z4/z1/_00_ ));
 sky130_fd_sc_hd__conb_1 \v0/z4/z1/_12_  (.LO(\v0/z4/z1/_01_ ));
 sky130_fd_sc_hd__conb_1 \v0/z4/z1/_13_  (.LO(\v0/z4/z1/_02_ ));
 sky130_fd_sc_hd__conb_1 \v0/z4/z1/_14_  (.LO(\v0/z4/z1/_03_ ));
 sky130_fd_sc_hd__conb_1 \v0/z4/z1/_15_  (.LO(\v0/z4/z1/_04_ ));
 sky130_fd_sc_hd__conb_1 \v0/z4/z1/_16_  (.LO(\v0/z4/z1/_05_ ));
 sky130_fd_sc_hd__conb_1 \v0/z4/z1/_17_  (.LO(\v0/z4/z1/_06_ ));
 sky130_fd_sc_hd__conb_1 \v0/z4/z1/_18_  (.LO(\v0/z4/z1/_07_ ));
 sky130_fd_sc_hd__conb_1 \v0/z4/z1/_19_  (.LO(\v0/z4/z1/_08_ ));
 sky130_fd_sc_hd__conb_1 \v0/z4/z1/_20_  (.LO(\v0/z4/z1/_09_ ));
 sky130_fd_sc_hd__conb_1 \v0/z4/z1/_21_  (.LO(\v0/z4/z1/_10_ ));
 sky130_fd_sc_hd__and2_0 \v0/z4/z1/z1/_0_  (.A(abs_b[8]),
    .B(abs_a[8]),
    .X(\v0/q3 [0]));
 sky130_fd_sc_hd__and2_0 \v0/z4/z1/z1/_1_  (.A(abs_b[8]),
    .B(abs_a[9]),
    .X(\v0/z4/z1/z1/temp [0]));
 sky130_fd_sc_hd__and2_0 \v0/z4/z1/z1/_2_  (.A(abs_a[8]),
    .B(abs_b[9]),
    .X(\v0/z4/z1/z1/temp [1]));
 sky130_fd_sc_hd__and2_0 \v0/z4/z1/z1/_3_  (.A(abs_a[9]),
    .B(abs_b[9]),
    .X(\v0/z4/z1/z1/temp [2]));
 sky130_fd_sc_hd__and2_0 \v0/z4/z1/z1/z1/_0_  (.A(\v0/z4/z1/z1/temp [1]),
    .B(\v0/z4/z1/z1/temp [0]),
    .X(\v0/z4/z1/z1/temp [3]));
 sky130_fd_sc_hd__xor2_1 \v0/z4/z1/z1/z1/_1_  (.A(\v0/z4/z1/z1/temp [1]),
    .B(\v0/z4/z1/z1/temp [0]),
    .X(\v0/q3 [1]));
 sky130_fd_sc_hd__and2_0 \v0/z4/z1/z1/z2/_0_  (.A(\v0/z4/z1/z1/temp [3]),
    .B(\v0/z4/z1/z1/temp [2]),
    .X(\v0/z4/z1/q0 [3]));
 sky130_fd_sc_hd__xor2_1 \v0/z4/z1/z1/z2/_1_  (.A(\v0/z4/z1/z1/temp [3]),
    .B(\v0/z4/z1/z1/temp [2]),
    .X(\v0/z4/z1/q0 [2]));
 sky130_fd_sc_hd__and2_0 \v0/z4/z1/z2/_0_  (.A(abs_b[8]),
    .B(abs_a[10]),
    .X(\v0/z4/z1/q1 [0]));
 sky130_fd_sc_hd__and2_0 \v0/z4/z1/z2/_1_  (.A(abs_b[8]),
    .B(abs_a[11]),
    .X(\v0/z4/z1/z2/temp [0]));
 sky130_fd_sc_hd__and2_0 \v0/z4/z1/z2/_2_  (.A(abs_a[10]),
    .B(abs_b[9]),
    .X(\v0/z4/z1/z2/temp [1]));
 sky130_fd_sc_hd__and2_0 \v0/z4/z1/z2/_3_  (.A(abs_a[11]),
    .B(abs_b[9]),
    .X(\v0/z4/z1/z2/temp [2]));
 sky130_fd_sc_hd__and2_0 \v0/z4/z1/z2/z1/_0_  (.A(\v0/z4/z1/z2/temp [1]),
    .B(\v0/z4/z1/z2/temp [0]),
    .X(\v0/z4/z1/z2/temp [3]));
 sky130_fd_sc_hd__xor2_1 \v0/z4/z1/z2/z1/_1_  (.A(\v0/z4/z1/z2/temp [1]),
    .B(\v0/z4/z1/z2/temp [0]),
    .X(\v0/z4/z1/q1 [1]));
 sky130_fd_sc_hd__and2_0 \v0/z4/z1/z2/z2/_0_  (.A(\v0/z4/z1/z2/temp [3]),
    .B(\v0/z4/z1/z2/temp [2]),
    .X(\v0/z4/z1/q1 [3]));
 sky130_fd_sc_hd__xor2_1 \v0/z4/z1/z2/z2/_1_  (.A(\v0/z4/z1/z2/temp [3]),
    .B(\v0/z4/z1/z2/temp [2]),
    .X(\v0/z4/z1/q1 [2]));
 sky130_fd_sc_hd__and2_0 \v0/z4/z1/z3/_0_  (.A(abs_b[10]),
    .B(abs_a[8]),
    .X(\v0/z4/z1/q2 [0]));
 sky130_fd_sc_hd__and2_0 \v0/z4/z1/z3/_1_  (.A(abs_b[10]),
    .B(abs_a[9]),
    .X(\v0/z4/z1/z3/temp [0]));
 sky130_fd_sc_hd__and2_0 \v0/z4/z1/z3/_2_  (.A(abs_a[8]),
    .B(abs_b[11]),
    .X(\v0/z4/z1/z3/temp [1]));
 sky130_fd_sc_hd__and2_0 \v0/z4/z1/z3/_3_  (.A(abs_a[9]),
    .B(abs_b[11]),
    .X(\v0/z4/z1/z3/temp [2]));
 sky130_fd_sc_hd__and2_0 \v0/z4/z1/z3/z1/_0_  (.A(\v0/z4/z1/z3/temp [1]),
    .B(\v0/z4/z1/z3/temp [0]),
    .X(\v0/z4/z1/z3/temp [3]));
 sky130_fd_sc_hd__xor2_1 \v0/z4/z1/z3/z1/_1_  (.A(\v0/z4/z1/z3/temp [1]),
    .B(\v0/z4/z1/z3/temp [0]),
    .X(\v0/z4/z1/q2 [1]));
 sky130_fd_sc_hd__and2_0 \v0/z4/z1/z3/z2/_0_  (.A(\v0/z4/z1/z3/temp [3]),
    .B(\v0/z4/z1/z3/temp [2]),
    .X(\v0/z4/z1/q2 [3]));
 sky130_fd_sc_hd__xor2_1 \v0/z4/z1/z3/z2/_1_  (.A(\v0/z4/z1/z3/temp [3]),
    .B(\v0/z4/z1/z3/temp [2]),
    .X(\v0/z4/z1/q2 [2]));
 sky130_fd_sc_hd__and2_0 \v0/z4/z1/z4/_0_  (.A(abs_b[10]),
    .B(abs_a[10]),
    .X(\v0/z4/z1/q3 [0]));
 sky130_fd_sc_hd__and2_0 \v0/z4/z1/z4/_1_  (.A(abs_b[10]),
    .B(abs_a[11]),
    .X(\v0/z4/z1/z4/temp [0]));
 sky130_fd_sc_hd__and2_0 \v0/z4/z1/z4/_2_  (.A(abs_a[10]),
    .B(abs_b[11]),
    .X(\v0/z4/z1/z4/temp [1]));
 sky130_fd_sc_hd__and2_0 \v0/z4/z1/z4/_3_  (.A(abs_a[11]),
    .B(abs_b[11]),
    .X(\v0/z4/z1/z4/temp [2]));
 sky130_fd_sc_hd__and2_0 \v0/z4/z1/z4/z1/_0_  (.A(\v0/z4/z1/z4/temp [1]),
    .B(\v0/z4/z1/z4/temp [0]),
    .X(\v0/z4/z1/z4/temp [3]));
 sky130_fd_sc_hd__xor2_1 \v0/z4/z1/z4/z1/_1_  (.A(\v0/z4/z1/z4/temp [1]),
    .B(\v0/z4/z1/z4/temp [0]),
    .X(\v0/z4/z1/q3 [1]));
 sky130_fd_sc_hd__and2_0 \v0/z4/z1/z4/z2/_0_  (.A(\v0/z4/z1/z4/temp [3]),
    .B(\v0/z4/z1/z4/temp [2]),
    .X(\v0/z4/z1/q3 [3]));
 sky130_fd_sc_hd__xor2_1 \v0/z4/z1/z4/z2/_1_  (.A(\v0/z4/z1/z4/temp [3]),
    .B(\v0/z4/z1/z4/temp [2]),
    .X(\v0/z4/z1/q3 [2]));
 sky130_fd_sc_hd__xnor2_1 \v0/z4/z1/z5/_07_  (.A(\v0/z4/z1/q0 [2]),
    .B(\v0/z4/z1/q1 [0]),
    .Y(\v0/z4/z1/z5/_00_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z4/z1/z5/_08_  (.A(\v0/z4/z1/_02_ ),
    .B(\v0/z4/z1/z5/_00_ ),
    .Y(\v0/z4/z1/q4 [0]));
 sky130_fd_sc_hd__maj3_1 \v0/z4/z1/z5/_09_  (.A(\v0/z4/z1/q0 [2]),
    .B(\v0/z4/z1/q1 [0]),
    .C(\v0/z4/z1/_02_ ),
    .X(\v0/z4/z1/z5/_01_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z4/z1/z5/_10_  (.A(\v0/z4/z1/q0 [3]),
    .B(\v0/z4/z1/q1 [1]),
    .Y(\v0/z4/z1/z5/_02_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z4/z1/z5/_11_  (.A(\v0/z4/z1/z5/_01_ ),
    .B(\v0/z4/z1/z5/_02_ ),
    .Y(\v0/z4/z1/q4 [1]));
 sky130_fd_sc_hd__maj3_1 \v0/z4/z1/z5/_12_  (.A(\v0/z4/z1/q0 [3]),
    .B(\v0/z4/z1/q1 [1]),
    .C(\v0/z4/z1/z5/_01_ ),
    .X(\v0/z4/z1/z5/_03_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z4/z1/z5/_13_  (.A(\v0/z4/z1/_00_ ),
    .B(\v0/z4/z1/q1 [2]),
    .Y(\v0/z4/z1/z5/_04_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z4/z1/z5/_14_  (.A(\v0/z4/z1/z5/_03_ ),
    .B(\v0/z4/z1/z5/_04_ ),
    .Y(\v0/z4/z1/q4 [2]));
 sky130_fd_sc_hd__maj3_1 \v0/z4/z1/z5/_15_  (.A(\v0/z4/z1/_00_ ),
    .B(\v0/z4/z1/q1 [2]),
    .C(\v0/z4/z1/z5/_03_ ),
    .X(\v0/z4/z1/z5/_05_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z4/z1/z5/_16_  (.A(\v0/z4/z1/_01_ ),
    .B(\v0/z4/z1/q1 [3]),
    .Y(\v0/z4/z1/z5/_06_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z4/z1/z5/_17_  (.A(\v0/z4/z1/z5/_05_ ),
    .B(\v0/z4/z1/z5/_06_ ),
    .Y(\v0/z4/z1/q4 [3]));
 sky130_fd_sc_hd__maj3_1 \v0/z4/z1/z5/_18_  (.A(\v0/z4/z1/_01_ ),
    .B(\v0/z4/z1/q1 [3]),
    .C(\v0/z4/z1/z5/_05_ ),
    .X(\v0/z4/z1/z5/Cout ));
 sky130_fd_sc_hd__xnor2_1 \v0/z4/z1/z6/_19_  (.A(\v0/z4/z1/_05_ ),
    .B(\v0/z4/z1/q2 [0]),
    .Y(\v0/z4/z1/z6/_00_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z4/z1/z6/_20_  (.A(\v0/z4/z1/_07_ ),
    .B(\v0/z4/z1/z6/_00_ ),
    .Y(\v0/z4/z1/q5 [0]));
 sky130_fd_sc_hd__maj3_1 \v0/z4/z1/z6/_21_  (.A(\v0/z4/z1/_05_ ),
    .B(\v0/z4/z1/q2 [0]),
    .C(\v0/z4/z1/_07_ ),
    .X(\v0/z4/z1/z6/_01_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z4/z1/z6/_22_  (.A(\v0/z4/z1/_06_ ),
    .B(\v0/z4/z1/q2 [1]),
    .Y(\v0/z4/z1/z6/_02_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z4/z1/z6/_23_  (.A(\v0/z4/z1/z6/_01_ ),
    .B(\v0/z4/z1/z6/_02_ ),
    .Y(\v0/z4/z1/q5 [1]));
 sky130_fd_sc_hd__maj3_1 \v0/z4/z1/z6/_24_  (.A(\v0/z4/z1/_06_ ),
    .B(\v0/z4/z1/q2 [1]),
    .C(\v0/z4/z1/z6/_01_ ),
    .X(\v0/z4/z1/z6/_03_ ));
 sky130_fd_sc_hd__lpflow_inputiso1p_1 \v0/z4/z1/z6/_25_  (.A(\v0/z4/z1/q3 [0]),
    .SLEEP(\v0/z4/z1/q2 [2]),
    .X(\v0/z4/z1/z6/_04_ ));
 sky130_fd_sc_hd__and2_0 \v0/z4/z1/z6/_26_  (.A(\v0/z4/z1/q3 [0]),
    .B(\v0/z4/z1/q2 [2]),
    .X(\v0/z4/z1/z6/_05_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z4/z1/z6/_27_  (.A(\v0/z4/z1/q3 [0]),
    .B(\v0/z4/z1/q2 [2]),
    .Y(\v0/z4/z1/z6/_06_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z4/z1/z6/_28_  (.A(\v0/z4/z1/z6/_04_ ),
    .B(\v0/z4/z1/z6/_06_ ),
    .Y(\v0/z4/z1/z6/_07_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z4/z1/z6/_29_  (.A(\v0/z4/z1/z6/_03_ ),
    .B(\v0/z4/z1/z6/_07_ ),
    .Y(\v0/z4/z1/q5 [2]));
 sky130_fd_sc_hd__nand2_1 \v0/z4/z1/z6/_30_  (.A(\v0/z4/z1/q3 [1]),
    .B(\v0/z4/z1/q2 [3]),
    .Y(\v0/z4/z1/z6/_08_ ));
 sky130_fd_sc_hd__xor2_1 \v0/z4/z1/z6/_31_  (.A(\v0/z4/z1/q3 [1]),
    .B(\v0/z4/z1/q2 [3]),
    .X(\v0/z4/z1/z6/_09_ ));
 sky130_fd_sc_hd__o21ai_0 \v0/z4/z1/z6/_32_  (.A1(\v0/z4/z1/z6/_03_ ),
    .A2(\v0/z4/z1/z6/_05_ ),
    .B1(\v0/z4/z1/z6/_04_ ),
    .Y(\v0/z4/z1/z6/_10_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z4/z1/z6/_33_  (.A(\v0/z4/z1/z6/_09_ ),
    .B(\v0/z4/z1/z6/_10_ ),
    .Y(\v0/z4/z1/q5 [3]));
 sky130_fd_sc_hd__nor2_1 \v0/z4/z1/z6/_34_  (.A(\v0/z4/z1/q3 [2]),
    .B(\v0/z4/z1/_03_ ),
    .Y(\v0/z4/z1/z6/_11_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z4/z1/z6/_35_  (.A(\v0/z4/z1/q3 [2]),
    .B(\v0/z4/z1/_03_ ),
    .Y(\v0/z4/z1/z6/_12_ ));
 sky130_fd_sc_hd__nand2b_1 \v0/z4/z1/z6/_36_  (.A_N(\v0/z4/z1/z6/_11_ ),
    .B(\v0/z4/z1/z6/_12_ ),
    .Y(\v0/z4/z1/z6/_13_ ));
 sky130_fd_sc_hd__o221ai_1 \v0/z4/z1/z6/_37_  (.A1(\v0/z4/z1/q3 [1]),
    .A2(\v0/z4/z1/q2 [3]),
    .B1(\v0/z4/z1/z6/_03_ ),
    .B2(\v0/z4/z1/z6/_05_ ),
    .C1(\v0/z4/z1/z6/_04_ ),
    .Y(\v0/z4/z1/z6/_14_ ));
 sky130_fd_sc_hd__a21oi_1 \v0/z4/z1/z6/_38_  (.A1(\v0/z4/z1/z6/_08_ ),
    .A2(\v0/z4/z1/z6/_14_ ),
    .B1(\v0/z4/z1/z6/_13_ ),
    .Y(\v0/z4/z1/z6/_15_ ));
 sky130_fd_sc_hd__and3_1 \v0/z4/z1/z6/_39_  (.A(\v0/z4/z1/z6/_08_ ),
    .B(\v0/z4/z1/z6/_13_ ),
    .C(\v0/z4/z1/z6/_14_ ),
    .X(\v0/z4/z1/z6/_16_ ));
 sky130_fd_sc_hd__nor2_1 \v0/z4/z1/z6/_40_  (.A(\v0/z4/z1/z6/_15_ ),
    .B(\v0/z4/z1/z6/_16_ ),
    .Y(\v0/z4/z1/q5 [4]));
 sky130_fd_sc_hd__xnor2_1 \v0/z4/z1/z6/_41_  (.A(\v0/z4/z1/q3 [3]),
    .B(\v0/z4/z1/_04_ ),
    .Y(\v0/z4/z1/z6/_17_ ));
 sky130_fd_sc_hd__a31oi_1 \v0/z4/z1/z6/_42_  (.A1(\v0/z4/z1/z6/_08_ ),
    .A2(\v0/z4/z1/z6/_12_ ),
    .A3(\v0/z4/z1/z6/_14_ ),
    .B1(\v0/z4/z1/z6/_11_ ),
    .Y(\v0/z4/z1/z6/_18_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z4/z1/z6/_43_  (.A(\v0/z4/z1/z6/_17_ ),
    .B(\v0/z4/z1/z6/_18_ ),
    .Y(\v0/z4/z1/q5 [5]));
 sky130_fd_sc_hd__maj3_1 \v0/z4/z1/z6/_44_  (.A(\v0/z4/z1/q3 [3]),
    .B(\v0/z4/z1/_04_ ),
    .C(\v0/z4/z1/z6/_18_ ),
    .X(\v0/z4/z1/z6/Cout ));
 sky130_fd_sc_hd__xnor2_1 \v0/z4/z1/z7/_19_  (.A(\v0/z4/z1/q5 [0]),
    .B(\v0/z4/z1/q4 [0]),
    .Y(\v0/z4/z1/z7/_00_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z4/z1/z7/_20_  (.A(\v0/z4/z1/_10_ ),
    .B(\v0/z4/z1/z7/_00_ ),
    .Y(\v0/q3 [2]));
 sky130_fd_sc_hd__maj3_1 \v0/z4/z1/z7/_21_  (.A(\v0/z4/z1/q5 [0]),
    .B(\v0/z4/z1/q4 [0]),
    .C(\v0/z4/z1/_10_ ),
    .X(\v0/z4/z1/z7/_01_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z4/z1/z7/_22_  (.A(\v0/z4/z1/q5 [1]),
    .B(\v0/z4/z1/q4 [1]),
    .Y(\v0/z4/z1/z7/_02_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z4/z1/z7/_23_  (.A(\v0/z4/z1/z7/_01_ ),
    .B(\v0/z4/z1/z7/_02_ ),
    .Y(\v0/q3 [3]));
 sky130_fd_sc_hd__maj3_1 \v0/z4/z1/z7/_24_  (.A(\v0/z4/z1/q5 [1]),
    .B(\v0/z4/z1/q4 [1]),
    .C(\v0/z4/z1/z7/_01_ ),
    .X(\v0/z4/z1/z7/_03_ ));
 sky130_fd_sc_hd__lpflow_inputiso1p_1 \v0/z4/z1/z7/_25_  (.A(\v0/z4/z1/q5 [2]),
    .SLEEP(\v0/z4/z1/q4 [2]),
    .X(\v0/z4/z1/z7/_04_ ));
 sky130_fd_sc_hd__and2_0 \v0/z4/z1/z7/_26_  (.A(\v0/z4/z1/q5 [2]),
    .B(\v0/z4/z1/q4 [2]),
    .X(\v0/z4/z1/z7/_05_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z4/z1/z7/_27_  (.A(\v0/z4/z1/q5 [2]),
    .B(\v0/z4/z1/q4 [2]),
    .Y(\v0/z4/z1/z7/_06_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z4/z1/z7/_28_  (.A(\v0/z4/z1/z7/_04_ ),
    .B(\v0/z4/z1/z7/_06_ ),
    .Y(\v0/z4/z1/z7/_07_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z4/z1/z7/_29_  (.A(\v0/z4/z1/z7/_03_ ),
    .B(\v0/z4/z1/z7/_07_ ),
    .Y(\v0/z4/q0 [4]));
 sky130_fd_sc_hd__nand2_1 \v0/z4/z1/z7/_30_  (.A(\v0/z4/z1/q5 [3]),
    .B(\v0/z4/z1/q4 [3]),
    .Y(\v0/z4/z1/z7/_08_ ));
 sky130_fd_sc_hd__xor2_1 \v0/z4/z1/z7/_31_  (.A(\v0/z4/z1/q5 [3]),
    .B(\v0/z4/z1/q4 [3]),
    .X(\v0/z4/z1/z7/_09_ ));
 sky130_fd_sc_hd__o21ai_0 \v0/z4/z1/z7/_32_  (.A1(\v0/z4/z1/z7/_03_ ),
    .A2(\v0/z4/z1/z7/_05_ ),
    .B1(\v0/z4/z1/z7/_04_ ),
    .Y(\v0/z4/z1/z7/_10_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z4/z1/z7/_33_  (.A(\v0/z4/z1/z7/_09_ ),
    .B(\v0/z4/z1/z7/_10_ ),
    .Y(\v0/z4/q0 [5]));
 sky130_fd_sc_hd__nor2_1 \v0/z4/z1/z7/_34_  (.A(\v0/z4/z1/q5 [4]),
    .B(\v0/z4/z1/_08_ ),
    .Y(\v0/z4/z1/z7/_11_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z4/z1/z7/_35_  (.A(\v0/z4/z1/q5 [4]),
    .B(\v0/z4/z1/_08_ ),
    .Y(\v0/z4/z1/z7/_12_ ));
 sky130_fd_sc_hd__nand2b_1 \v0/z4/z1/z7/_36_  (.A_N(\v0/z4/z1/z7/_11_ ),
    .B(\v0/z4/z1/z7/_12_ ),
    .Y(\v0/z4/z1/z7/_13_ ));
 sky130_fd_sc_hd__o221ai_1 \v0/z4/z1/z7/_37_  (.A1(\v0/z4/z1/q5 [3]),
    .A2(\v0/z4/z1/q4 [3]),
    .B1(\v0/z4/z1/z7/_03_ ),
    .B2(\v0/z4/z1/z7/_05_ ),
    .C1(\v0/z4/z1/z7/_04_ ),
    .Y(\v0/z4/z1/z7/_14_ ));
 sky130_fd_sc_hd__a21oi_1 \v0/z4/z1/z7/_38_  (.A1(\v0/z4/z1/z7/_08_ ),
    .A2(\v0/z4/z1/z7/_14_ ),
    .B1(\v0/z4/z1/z7/_13_ ),
    .Y(\v0/z4/z1/z7/_15_ ));
 sky130_fd_sc_hd__and3_1 \v0/z4/z1/z7/_39_  (.A(\v0/z4/z1/z7/_08_ ),
    .B(\v0/z4/z1/z7/_13_ ),
    .C(\v0/z4/z1/z7/_14_ ),
    .X(\v0/z4/z1/z7/_16_ ));
 sky130_fd_sc_hd__nor2_1 \v0/z4/z1/z7/_40_  (.A(\v0/z4/z1/z7/_15_ ),
    .B(\v0/z4/z1/z7/_16_ ),
    .Y(\v0/z4/q0 [6]));
 sky130_fd_sc_hd__xnor2_1 \v0/z4/z1/z7/_41_  (.A(\v0/z4/z1/q5 [5]),
    .B(\v0/z4/z1/_09_ ),
    .Y(\v0/z4/z1/z7/_17_ ));
 sky130_fd_sc_hd__a31oi_1 \v0/z4/z1/z7/_42_  (.A1(\v0/z4/z1/z7/_08_ ),
    .A2(\v0/z4/z1/z7/_12_ ),
    .A3(\v0/z4/z1/z7/_14_ ),
    .B1(\v0/z4/z1/z7/_11_ ),
    .Y(\v0/z4/z1/z7/_18_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z4/z1/z7/_43_  (.A(\v0/z4/z1/z7/_17_ ),
    .B(\v0/z4/z1/z7/_18_ ),
    .Y(\v0/z4/q0 [7]));
 sky130_fd_sc_hd__maj3_1 \v0/z4/z1/z7/_44_  (.A(\v0/z4/z1/q5 [5]),
    .B(\v0/z4/z1/_09_ ),
    .C(\v0/z4/z1/z7/_18_ ),
    .X(\v0/z4/z1/z7/Cout ));
 sky130_fd_sc_hd__conb_1 \v0/z4/z2/_11_  (.LO(\v0/z4/z2/_00_ ));
 sky130_fd_sc_hd__conb_1 \v0/z4/z2/_12_  (.LO(\v0/z4/z2/_01_ ));
 sky130_fd_sc_hd__conb_1 \v0/z4/z2/_13_  (.LO(\v0/z4/z2/_02_ ));
 sky130_fd_sc_hd__conb_1 \v0/z4/z2/_14_  (.LO(\v0/z4/z2/_03_ ));
 sky130_fd_sc_hd__conb_1 \v0/z4/z2/_15_  (.LO(\v0/z4/z2/_04_ ));
 sky130_fd_sc_hd__conb_1 \v0/z4/z2/_16_  (.LO(\v0/z4/z2/_05_ ));
 sky130_fd_sc_hd__conb_1 \v0/z4/z2/_17_  (.LO(\v0/z4/z2/_06_ ));
 sky130_fd_sc_hd__conb_1 \v0/z4/z2/_18_  (.LO(\v0/z4/z2/_07_ ));
 sky130_fd_sc_hd__conb_1 \v0/z4/z2/_19_  (.LO(\v0/z4/z2/_08_ ));
 sky130_fd_sc_hd__conb_1 \v0/z4/z2/_20_  (.LO(\v0/z4/z2/_09_ ));
 sky130_fd_sc_hd__conb_1 \v0/z4/z2/_21_  (.LO(\v0/z4/z2/_10_ ));
 sky130_fd_sc_hd__and2_0 \v0/z4/z2/z1/_0_  (.A(abs_b[8]),
    .B(abs_a[12]),
    .X(\v0/z4/q1 [0]));
 sky130_fd_sc_hd__and2_0 \v0/z4/z2/z1/_1_  (.A(abs_b[8]),
    .B(abs_a[13]),
    .X(\v0/z4/z2/z1/temp [0]));
 sky130_fd_sc_hd__and2_0 \v0/z4/z2/z1/_2_  (.A(abs_a[12]),
    .B(abs_b[9]),
    .X(\v0/z4/z2/z1/temp [1]));
 sky130_fd_sc_hd__and2_0 \v0/z4/z2/z1/_3_  (.A(abs_a[13]),
    .B(abs_b[9]),
    .X(\v0/z4/z2/z1/temp [2]));
 sky130_fd_sc_hd__and2_0 \v0/z4/z2/z1/z1/_0_  (.A(\v0/z4/z2/z1/temp [1]),
    .B(\v0/z4/z2/z1/temp [0]),
    .X(\v0/z4/z2/z1/temp [3]));
 sky130_fd_sc_hd__xor2_1 \v0/z4/z2/z1/z1/_1_  (.A(\v0/z4/z2/z1/temp [1]),
    .B(\v0/z4/z2/z1/temp [0]),
    .X(\v0/z4/q1 [1]));
 sky130_fd_sc_hd__and2_0 \v0/z4/z2/z1/z2/_0_  (.A(\v0/z4/z2/z1/temp [3]),
    .B(\v0/z4/z2/z1/temp [2]),
    .X(\v0/z4/z2/q0 [3]));
 sky130_fd_sc_hd__xor2_1 \v0/z4/z2/z1/z2/_1_  (.A(\v0/z4/z2/z1/temp [3]),
    .B(\v0/z4/z2/z1/temp [2]),
    .X(\v0/z4/z2/q0 [2]));
 sky130_fd_sc_hd__and2_0 \v0/z4/z2/z2/_0_  (.A(abs_b[8]),
    .B(abs_a[14]),
    .X(\v0/z4/z2/q1 [0]));
 sky130_fd_sc_hd__and2_0 \v0/z4/z2/z2/_1_  (.A(abs_b[8]),
    .B(abs_a[15]),
    .X(\v0/z4/z2/z2/temp [0]));
 sky130_fd_sc_hd__and2_0 \v0/z4/z2/z2/_2_  (.A(abs_a[14]),
    .B(abs_b[9]),
    .X(\v0/z4/z2/z2/temp [1]));
 sky130_fd_sc_hd__and2_0 \v0/z4/z2/z2/_3_  (.A(abs_a[15]),
    .B(abs_b[9]),
    .X(\v0/z4/z2/z2/temp [2]));
 sky130_fd_sc_hd__and2_0 \v0/z4/z2/z2/z1/_0_  (.A(\v0/z4/z2/z2/temp [1]),
    .B(\v0/z4/z2/z2/temp [0]),
    .X(\v0/z4/z2/z2/temp [3]));
 sky130_fd_sc_hd__xor2_1 \v0/z4/z2/z2/z1/_1_  (.A(\v0/z4/z2/z2/temp [1]),
    .B(\v0/z4/z2/z2/temp [0]),
    .X(\v0/z4/z2/q1 [1]));
 sky130_fd_sc_hd__and2_0 \v0/z4/z2/z2/z2/_0_  (.A(\v0/z4/z2/z2/temp [3]),
    .B(\v0/z4/z2/z2/temp [2]),
    .X(\v0/z4/z2/q1 [3]));
 sky130_fd_sc_hd__xor2_1 \v0/z4/z2/z2/z2/_1_  (.A(\v0/z4/z2/z2/temp [3]),
    .B(\v0/z4/z2/z2/temp [2]),
    .X(\v0/z4/z2/q1 [2]));
 sky130_fd_sc_hd__and2_0 \v0/z4/z2/z3/_0_  (.A(abs_b[10]),
    .B(abs_a[12]),
    .X(\v0/z4/z2/q2 [0]));
 sky130_fd_sc_hd__and2_0 \v0/z4/z2/z3/_1_  (.A(abs_b[10]),
    .B(abs_a[13]),
    .X(\v0/z4/z2/z3/temp [0]));
 sky130_fd_sc_hd__and2_0 \v0/z4/z2/z3/_2_  (.A(abs_a[12]),
    .B(abs_b[11]),
    .X(\v0/z4/z2/z3/temp [1]));
 sky130_fd_sc_hd__and2_0 \v0/z4/z2/z3/_3_  (.A(abs_a[13]),
    .B(abs_b[11]),
    .X(\v0/z4/z2/z3/temp [2]));
 sky130_fd_sc_hd__and2_0 \v0/z4/z2/z3/z1/_0_  (.A(\v0/z4/z2/z3/temp [1]),
    .B(\v0/z4/z2/z3/temp [0]),
    .X(\v0/z4/z2/z3/temp [3]));
 sky130_fd_sc_hd__xor2_1 \v0/z4/z2/z3/z1/_1_  (.A(\v0/z4/z2/z3/temp [1]),
    .B(\v0/z4/z2/z3/temp [0]),
    .X(\v0/z4/z2/q2 [1]));
 sky130_fd_sc_hd__and2_0 \v0/z4/z2/z3/z2/_0_  (.A(\v0/z4/z2/z3/temp [3]),
    .B(\v0/z4/z2/z3/temp [2]),
    .X(\v0/z4/z2/q2 [3]));
 sky130_fd_sc_hd__xor2_1 \v0/z4/z2/z3/z2/_1_  (.A(\v0/z4/z2/z3/temp [3]),
    .B(\v0/z4/z2/z3/temp [2]),
    .X(\v0/z4/z2/q2 [2]));
 sky130_fd_sc_hd__and2_0 \v0/z4/z2/z4/_0_  (.A(abs_b[10]),
    .B(abs_a[14]),
    .X(\v0/z4/z2/q3 [0]));
 sky130_fd_sc_hd__and2_0 \v0/z4/z2/z4/_1_  (.A(abs_b[10]),
    .B(abs_a[15]),
    .X(\v0/z4/z2/z4/temp [0]));
 sky130_fd_sc_hd__and2_0 \v0/z4/z2/z4/_2_  (.A(abs_a[14]),
    .B(abs_b[11]),
    .X(\v0/z4/z2/z4/temp [1]));
 sky130_fd_sc_hd__and2_0 \v0/z4/z2/z4/_3_  (.A(abs_a[15]),
    .B(abs_b[11]),
    .X(\v0/z4/z2/z4/temp [2]));
 sky130_fd_sc_hd__and2_0 \v0/z4/z2/z4/z1/_0_  (.A(\v0/z4/z2/z4/temp [1]),
    .B(\v0/z4/z2/z4/temp [0]),
    .X(\v0/z4/z2/z4/temp [3]));
 sky130_fd_sc_hd__xor2_1 \v0/z4/z2/z4/z1/_1_  (.A(\v0/z4/z2/z4/temp [1]),
    .B(\v0/z4/z2/z4/temp [0]),
    .X(\v0/z4/z2/q3 [1]));
 sky130_fd_sc_hd__and2_0 \v0/z4/z2/z4/z2/_0_  (.A(\v0/z4/z2/z4/temp [3]),
    .B(\v0/z4/z2/z4/temp [2]),
    .X(\v0/z4/z2/q3 [3]));
 sky130_fd_sc_hd__xor2_1 \v0/z4/z2/z4/z2/_1_  (.A(\v0/z4/z2/z4/temp [3]),
    .B(\v0/z4/z2/z4/temp [2]),
    .X(\v0/z4/z2/q3 [2]));
 sky130_fd_sc_hd__xnor2_1 \v0/z4/z2/z5/_07_  (.A(\v0/z4/z2/q0 [2]),
    .B(\v0/z4/z2/q1 [0]),
    .Y(\v0/z4/z2/z5/_00_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z4/z2/z5/_08_  (.A(\v0/z4/z2/_02_ ),
    .B(\v0/z4/z2/z5/_00_ ),
    .Y(\v0/z4/z2/q4 [0]));
 sky130_fd_sc_hd__maj3_1 \v0/z4/z2/z5/_09_  (.A(\v0/z4/z2/q0 [2]),
    .B(\v0/z4/z2/q1 [0]),
    .C(\v0/z4/z2/_02_ ),
    .X(\v0/z4/z2/z5/_01_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z4/z2/z5/_10_  (.A(\v0/z4/z2/q0 [3]),
    .B(\v0/z4/z2/q1 [1]),
    .Y(\v0/z4/z2/z5/_02_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z4/z2/z5/_11_  (.A(\v0/z4/z2/z5/_01_ ),
    .B(\v0/z4/z2/z5/_02_ ),
    .Y(\v0/z4/z2/q4 [1]));
 sky130_fd_sc_hd__maj3_1 \v0/z4/z2/z5/_12_  (.A(\v0/z4/z2/q0 [3]),
    .B(\v0/z4/z2/q1 [1]),
    .C(\v0/z4/z2/z5/_01_ ),
    .X(\v0/z4/z2/z5/_03_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z4/z2/z5/_13_  (.A(\v0/z4/z2/_00_ ),
    .B(\v0/z4/z2/q1 [2]),
    .Y(\v0/z4/z2/z5/_04_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z4/z2/z5/_14_  (.A(\v0/z4/z2/z5/_03_ ),
    .B(\v0/z4/z2/z5/_04_ ),
    .Y(\v0/z4/z2/q4 [2]));
 sky130_fd_sc_hd__maj3_1 \v0/z4/z2/z5/_15_  (.A(\v0/z4/z2/_00_ ),
    .B(\v0/z4/z2/q1 [2]),
    .C(\v0/z4/z2/z5/_03_ ),
    .X(\v0/z4/z2/z5/_05_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z4/z2/z5/_16_  (.A(\v0/z4/z2/_01_ ),
    .B(\v0/z4/z2/q1 [3]),
    .Y(\v0/z4/z2/z5/_06_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z4/z2/z5/_17_  (.A(\v0/z4/z2/z5/_05_ ),
    .B(\v0/z4/z2/z5/_06_ ),
    .Y(\v0/z4/z2/q4 [3]));
 sky130_fd_sc_hd__maj3_1 \v0/z4/z2/z5/_18_  (.A(\v0/z4/z2/_01_ ),
    .B(\v0/z4/z2/q1 [3]),
    .C(\v0/z4/z2/z5/_05_ ),
    .X(\v0/z4/z2/z5/Cout ));
 sky130_fd_sc_hd__xnor2_1 \v0/z4/z2/z6/_19_  (.A(\v0/z4/z2/_05_ ),
    .B(\v0/z4/z2/q2 [0]),
    .Y(\v0/z4/z2/z6/_00_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z4/z2/z6/_20_  (.A(\v0/z4/z2/_07_ ),
    .B(\v0/z4/z2/z6/_00_ ),
    .Y(\v0/z4/z2/q5 [0]));
 sky130_fd_sc_hd__maj3_1 \v0/z4/z2/z6/_21_  (.A(\v0/z4/z2/_05_ ),
    .B(\v0/z4/z2/q2 [0]),
    .C(\v0/z4/z2/_07_ ),
    .X(\v0/z4/z2/z6/_01_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z4/z2/z6/_22_  (.A(\v0/z4/z2/_06_ ),
    .B(\v0/z4/z2/q2 [1]),
    .Y(\v0/z4/z2/z6/_02_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z4/z2/z6/_23_  (.A(\v0/z4/z2/z6/_01_ ),
    .B(\v0/z4/z2/z6/_02_ ),
    .Y(\v0/z4/z2/q5 [1]));
 sky130_fd_sc_hd__maj3_1 \v0/z4/z2/z6/_24_  (.A(\v0/z4/z2/_06_ ),
    .B(\v0/z4/z2/q2 [1]),
    .C(\v0/z4/z2/z6/_01_ ),
    .X(\v0/z4/z2/z6/_03_ ));
 sky130_fd_sc_hd__lpflow_inputiso1p_1 \v0/z4/z2/z6/_25_  (.A(\v0/z4/z2/q3 [0]),
    .SLEEP(\v0/z4/z2/q2 [2]),
    .X(\v0/z4/z2/z6/_04_ ));
 sky130_fd_sc_hd__and2_0 \v0/z4/z2/z6/_26_  (.A(\v0/z4/z2/q3 [0]),
    .B(\v0/z4/z2/q2 [2]),
    .X(\v0/z4/z2/z6/_05_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z4/z2/z6/_27_  (.A(\v0/z4/z2/q3 [0]),
    .B(\v0/z4/z2/q2 [2]),
    .Y(\v0/z4/z2/z6/_06_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z4/z2/z6/_28_  (.A(\v0/z4/z2/z6/_04_ ),
    .B(\v0/z4/z2/z6/_06_ ),
    .Y(\v0/z4/z2/z6/_07_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z4/z2/z6/_29_  (.A(\v0/z4/z2/z6/_03_ ),
    .B(\v0/z4/z2/z6/_07_ ),
    .Y(\v0/z4/z2/q5 [2]));
 sky130_fd_sc_hd__nand2_1 \v0/z4/z2/z6/_30_  (.A(\v0/z4/z2/q3 [1]),
    .B(\v0/z4/z2/q2 [3]),
    .Y(\v0/z4/z2/z6/_08_ ));
 sky130_fd_sc_hd__xor2_1 \v0/z4/z2/z6/_31_  (.A(\v0/z4/z2/q3 [1]),
    .B(\v0/z4/z2/q2 [3]),
    .X(\v0/z4/z2/z6/_09_ ));
 sky130_fd_sc_hd__o21ai_0 \v0/z4/z2/z6/_32_  (.A1(\v0/z4/z2/z6/_03_ ),
    .A2(\v0/z4/z2/z6/_05_ ),
    .B1(\v0/z4/z2/z6/_04_ ),
    .Y(\v0/z4/z2/z6/_10_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z4/z2/z6/_33_  (.A(\v0/z4/z2/z6/_09_ ),
    .B(\v0/z4/z2/z6/_10_ ),
    .Y(\v0/z4/z2/q5 [3]));
 sky130_fd_sc_hd__nor2_1 \v0/z4/z2/z6/_34_  (.A(\v0/z4/z2/q3 [2]),
    .B(\v0/z4/z2/_03_ ),
    .Y(\v0/z4/z2/z6/_11_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z4/z2/z6/_35_  (.A(\v0/z4/z2/q3 [2]),
    .B(\v0/z4/z2/_03_ ),
    .Y(\v0/z4/z2/z6/_12_ ));
 sky130_fd_sc_hd__nand2b_1 \v0/z4/z2/z6/_36_  (.A_N(\v0/z4/z2/z6/_11_ ),
    .B(\v0/z4/z2/z6/_12_ ),
    .Y(\v0/z4/z2/z6/_13_ ));
 sky130_fd_sc_hd__o221ai_1 \v0/z4/z2/z6/_37_  (.A1(\v0/z4/z2/q3 [1]),
    .A2(\v0/z4/z2/q2 [3]),
    .B1(\v0/z4/z2/z6/_03_ ),
    .B2(\v0/z4/z2/z6/_05_ ),
    .C1(\v0/z4/z2/z6/_04_ ),
    .Y(\v0/z4/z2/z6/_14_ ));
 sky130_fd_sc_hd__a21oi_1 \v0/z4/z2/z6/_38_  (.A1(\v0/z4/z2/z6/_08_ ),
    .A2(\v0/z4/z2/z6/_14_ ),
    .B1(\v0/z4/z2/z6/_13_ ),
    .Y(\v0/z4/z2/z6/_15_ ));
 sky130_fd_sc_hd__and3_1 \v0/z4/z2/z6/_39_  (.A(\v0/z4/z2/z6/_08_ ),
    .B(\v0/z4/z2/z6/_13_ ),
    .C(\v0/z4/z2/z6/_14_ ),
    .X(\v0/z4/z2/z6/_16_ ));
 sky130_fd_sc_hd__nor2_1 \v0/z4/z2/z6/_40_  (.A(\v0/z4/z2/z6/_15_ ),
    .B(\v0/z4/z2/z6/_16_ ),
    .Y(\v0/z4/z2/q5 [4]));
 sky130_fd_sc_hd__xnor2_1 \v0/z4/z2/z6/_41_  (.A(\v0/z4/z2/q3 [3]),
    .B(\v0/z4/z2/_04_ ),
    .Y(\v0/z4/z2/z6/_17_ ));
 sky130_fd_sc_hd__a31oi_1 \v0/z4/z2/z6/_42_  (.A1(\v0/z4/z2/z6/_08_ ),
    .A2(\v0/z4/z2/z6/_12_ ),
    .A3(\v0/z4/z2/z6/_14_ ),
    .B1(\v0/z4/z2/z6/_11_ ),
    .Y(\v0/z4/z2/z6/_18_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z4/z2/z6/_43_  (.A(\v0/z4/z2/z6/_17_ ),
    .B(\v0/z4/z2/z6/_18_ ),
    .Y(\v0/z4/z2/q5 [5]));
 sky130_fd_sc_hd__maj3_1 \v0/z4/z2/z6/_44_  (.A(\v0/z4/z2/q3 [3]),
    .B(\v0/z4/z2/_04_ ),
    .C(\v0/z4/z2/z6/_18_ ),
    .X(\v0/z4/z2/z6/Cout ));
 sky130_fd_sc_hd__xnor2_1 \v0/z4/z2/z7/_19_  (.A(\v0/z4/z2/q5 [0]),
    .B(\v0/z4/z2/q4 [0]),
    .Y(\v0/z4/z2/z7/_00_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z4/z2/z7/_20_  (.A(\v0/z4/z2/_10_ ),
    .B(\v0/z4/z2/z7/_00_ ),
    .Y(\v0/z4/q1 [2]));
 sky130_fd_sc_hd__maj3_1 \v0/z4/z2/z7/_21_  (.A(\v0/z4/z2/q5 [0]),
    .B(\v0/z4/z2/q4 [0]),
    .C(\v0/z4/z2/_10_ ),
    .X(\v0/z4/z2/z7/_01_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z4/z2/z7/_22_  (.A(\v0/z4/z2/q5 [1]),
    .B(\v0/z4/z2/q4 [1]),
    .Y(\v0/z4/z2/z7/_02_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z4/z2/z7/_23_  (.A(\v0/z4/z2/z7/_01_ ),
    .B(\v0/z4/z2/z7/_02_ ),
    .Y(\v0/z4/q1 [3]));
 sky130_fd_sc_hd__maj3_1 \v0/z4/z2/z7/_24_  (.A(\v0/z4/z2/q5 [1]),
    .B(\v0/z4/z2/q4 [1]),
    .C(\v0/z4/z2/z7/_01_ ),
    .X(\v0/z4/z2/z7/_03_ ));
 sky130_fd_sc_hd__lpflow_inputiso1p_1 \v0/z4/z2/z7/_25_  (.A(\v0/z4/z2/q5 [2]),
    .SLEEP(\v0/z4/z2/q4 [2]),
    .X(\v0/z4/z2/z7/_04_ ));
 sky130_fd_sc_hd__and2_0 \v0/z4/z2/z7/_26_  (.A(\v0/z4/z2/q5 [2]),
    .B(\v0/z4/z2/q4 [2]),
    .X(\v0/z4/z2/z7/_05_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z4/z2/z7/_27_  (.A(\v0/z4/z2/q5 [2]),
    .B(\v0/z4/z2/q4 [2]),
    .Y(\v0/z4/z2/z7/_06_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z4/z2/z7/_28_  (.A(\v0/z4/z2/z7/_04_ ),
    .B(\v0/z4/z2/z7/_06_ ),
    .Y(\v0/z4/z2/z7/_07_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z4/z2/z7/_29_  (.A(\v0/z4/z2/z7/_03_ ),
    .B(\v0/z4/z2/z7/_07_ ),
    .Y(\v0/z4/q1 [4]));
 sky130_fd_sc_hd__nand2_1 \v0/z4/z2/z7/_30_  (.A(\v0/z4/z2/q5 [3]),
    .B(\v0/z4/z2/q4 [3]),
    .Y(\v0/z4/z2/z7/_08_ ));
 sky130_fd_sc_hd__xor2_1 \v0/z4/z2/z7/_31_  (.A(\v0/z4/z2/q5 [3]),
    .B(\v0/z4/z2/q4 [3]),
    .X(\v0/z4/z2/z7/_09_ ));
 sky130_fd_sc_hd__o21ai_0 \v0/z4/z2/z7/_32_  (.A1(\v0/z4/z2/z7/_03_ ),
    .A2(\v0/z4/z2/z7/_05_ ),
    .B1(\v0/z4/z2/z7/_04_ ),
    .Y(\v0/z4/z2/z7/_10_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z4/z2/z7/_33_  (.A(\v0/z4/z2/z7/_09_ ),
    .B(\v0/z4/z2/z7/_10_ ),
    .Y(\v0/z4/q1 [5]));
 sky130_fd_sc_hd__nor2_1 \v0/z4/z2/z7/_34_  (.A(\v0/z4/z2/q5 [4]),
    .B(\v0/z4/z2/_08_ ),
    .Y(\v0/z4/z2/z7/_11_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z4/z2/z7/_35_  (.A(\v0/z4/z2/q5 [4]),
    .B(\v0/z4/z2/_08_ ),
    .Y(\v0/z4/z2/z7/_12_ ));
 sky130_fd_sc_hd__nand2b_1 \v0/z4/z2/z7/_36_  (.A_N(\v0/z4/z2/z7/_11_ ),
    .B(\v0/z4/z2/z7/_12_ ),
    .Y(\v0/z4/z2/z7/_13_ ));
 sky130_fd_sc_hd__o221ai_1 \v0/z4/z2/z7/_37_  (.A1(\v0/z4/z2/q5 [3]),
    .A2(\v0/z4/z2/q4 [3]),
    .B1(\v0/z4/z2/z7/_03_ ),
    .B2(\v0/z4/z2/z7/_05_ ),
    .C1(\v0/z4/z2/z7/_04_ ),
    .Y(\v0/z4/z2/z7/_14_ ));
 sky130_fd_sc_hd__a21oi_1 \v0/z4/z2/z7/_38_  (.A1(\v0/z4/z2/z7/_08_ ),
    .A2(\v0/z4/z2/z7/_14_ ),
    .B1(\v0/z4/z2/z7/_13_ ),
    .Y(\v0/z4/z2/z7/_15_ ));
 sky130_fd_sc_hd__and3_1 \v0/z4/z2/z7/_39_  (.A(\v0/z4/z2/z7/_08_ ),
    .B(\v0/z4/z2/z7/_13_ ),
    .C(\v0/z4/z2/z7/_14_ ),
    .X(\v0/z4/z2/z7/_16_ ));
 sky130_fd_sc_hd__nor2_1 \v0/z4/z2/z7/_40_  (.A(\v0/z4/z2/z7/_15_ ),
    .B(\v0/z4/z2/z7/_16_ ),
    .Y(\v0/z4/q1 [6]));
 sky130_fd_sc_hd__xnor2_1 \v0/z4/z2/z7/_41_  (.A(\v0/z4/z2/q5 [5]),
    .B(\v0/z4/z2/_09_ ),
    .Y(\v0/z4/z2/z7/_17_ ));
 sky130_fd_sc_hd__a31oi_1 \v0/z4/z2/z7/_42_  (.A1(\v0/z4/z2/z7/_08_ ),
    .A2(\v0/z4/z2/z7/_12_ ),
    .A3(\v0/z4/z2/z7/_14_ ),
    .B1(\v0/z4/z2/z7/_11_ ),
    .Y(\v0/z4/z2/z7/_18_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z4/z2/z7/_43_  (.A(\v0/z4/z2/z7/_17_ ),
    .B(\v0/z4/z2/z7/_18_ ),
    .Y(\v0/z4/q1 [7]));
 sky130_fd_sc_hd__maj3_1 \v0/z4/z2/z7/_44_  (.A(\v0/z4/z2/q5 [5]),
    .B(\v0/z4/z2/_09_ ),
    .C(\v0/z4/z2/z7/_18_ ),
    .X(\v0/z4/z2/z7/Cout ));
 sky130_fd_sc_hd__conb_1 \v0/z4/z3/_11_  (.LO(\v0/z4/z3/_00_ ));
 sky130_fd_sc_hd__conb_1 \v0/z4/z3/_12_  (.LO(\v0/z4/z3/_01_ ));
 sky130_fd_sc_hd__conb_1 \v0/z4/z3/_13_  (.LO(\v0/z4/z3/_02_ ));
 sky130_fd_sc_hd__conb_1 \v0/z4/z3/_14_  (.LO(\v0/z4/z3/_03_ ));
 sky130_fd_sc_hd__conb_1 \v0/z4/z3/_15_  (.LO(\v0/z4/z3/_04_ ));
 sky130_fd_sc_hd__conb_1 \v0/z4/z3/_16_  (.LO(\v0/z4/z3/_05_ ));
 sky130_fd_sc_hd__conb_1 \v0/z4/z3/_17_  (.LO(\v0/z4/z3/_06_ ));
 sky130_fd_sc_hd__conb_1 \v0/z4/z3/_18_  (.LO(\v0/z4/z3/_07_ ));
 sky130_fd_sc_hd__conb_1 \v0/z4/z3/_19_  (.LO(\v0/z4/z3/_08_ ));
 sky130_fd_sc_hd__conb_1 \v0/z4/z3/_20_  (.LO(\v0/z4/z3/_09_ ));
 sky130_fd_sc_hd__conb_1 \v0/z4/z3/_21_  (.LO(\v0/z4/z3/_10_ ));
 sky130_fd_sc_hd__and2_0 \v0/z4/z3/z1/_0_  (.A(abs_b[12]),
    .B(abs_a[8]),
    .X(\v0/z4/q2 [0]));
 sky130_fd_sc_hd__and2_0 \v0/z4/z3/z1/_1_  (.A(abs_b[12]),
    .B(abs_a[9]),
    .X(\v0/z4/z3/z1/temp [0]));
 sky130_fd_sc_hd__and2_0 \v0/z4/z3/z1/_2_  (.A(abs_a[8]),
    .B(abs_b[13]),
    .X(\v0/z4/z3/z1/temp [1]));
 sky130_fd_sc_hd__and2_0 \v0/z4/z3/z1/_3_  (.A(abs_a[9]),
    .B(abs_b[13]),
    .X(\v0/z4/z3/z1/temp [2]));
 sky130_fd_sc_hd__and2_0 \v0/z4/z3/z1/z1/_0_  (.A(\v0/z4/z3/z1/temp [1]),
    .B(\v0/z4/z3/z1/temp [0]),
    .X(\v0/z4/z3/z1/temp [3]));
 sky130_fd_sc_hd__xor2_1 \v0/z4/z3/z1/z1/_1_  (.A(\v0/z4/z3/z1/temp [1]),
    .B(\v0/z4/z3/z1/temp [0]),
    .X(\v0/z4/q2 [1]));
 sky130_fd_sc_hd__and2_0 \v0/z4/z3/z1/z2/_0_  (.A(\v0/z4/z3/z1/temp [3]),
    .B(\v0/z4/z3/z1/temp [2]),
    .X(\v0/z4/z3/q0 [3]));
 sky130_fd_sc_hd__xor2_1 \v0/z4/z3/z1/z2/_1_  (.A(\v0/z4/z3/z1/temp [3]),
    .B(\v0/z4/z3/z1/temp [2]),
    .X(\v0/z4/z3/q0 [2]));
 sky130_fd_sc_hd__and2_0 \v0/z4/z3/z2/_0_  (.A(abs_b[12]),
    .B(abs_a[10]),
    .X(\v0/z4/z3/q1 [0]));
 sky130_fd_sc_hd__and2_0 \v0/z4/z3/z2/_1_  (.A(abs_b[12]),
    .B(abs_a[11]),
    .X(\v0/z4/z3/z2/temp [0]));
 sky130_fd_sc_hd__and2_0 \v0/z4/z3/z2/_2_  (.A(abs_a[10]),
    .B(abs_b[13]),
    .X(\v0/z4/z3/z2/temp [1]));
 sky130_fd_sc_hd__and2_0 \v0/z4/z3/z2/_3_  (.A(abs_a[11]),
    .B(abs_b[13]),
    .X(\v0/z4/z3/z2/temp [2]));
 sky130_fd_sc_hd__and2_0 \v0/z4/z3/z2/z1/_0_  (.A(\v0/z4/z3/z2/temp [1]),
    .B(\v0/z4/z3/z2/temp [0]),
    .X(\v0/z4/z3/z2/temp [3]));
 sky130_fd_sc_hd__xor2_1 \v0/z4/z3/z2/z1/_1_  (.A(\v0/z4/z3/z2/temp [1]),
    .B(\v0/z4/z3/z2/temp [0]),
    .X(\v0/z4/z3/q1 [1]));
 sky130_fd_sc_hd__and2_0 \v0/z4/z3/z2/z2/_0_  (.A(\v0/z4/z3/z2/temp [3]),
    .B(\v0/z4/z3/z2/temp [2]),
    .X(\v0/z4/z3/q1 [3]));
 sky130_fd_sc_hd__xor2_1 \v0/z4/z3/z2/z2/_1_  (.A(\v0/z4/z3/z2/temp [3]),
    .B(\v0/z4/z3/z2/temp [2]),
    .X(\v0/z4/z3/q1 [2]));
 sky130_fd_sc_hd__and2_0 \v0/z4/z3/z3/_0_  (.A(abs_b[14]),
    .B(abs_a[8]),
    .X(\v0/z4/z3/q2 [0]));
 sky130_fd_sc_hd__and2_0 \v0/z4/z3/z3/_1_  (.A(abs_b[14]),
    .B(abs_a[9]),
    .X(\v0/z4/z3/z3/temp [0]));
 sky130_fd_sc_hd__and2_0 \v0/z4/z3/z3/_2_  (.A(abs_a[8]),
    .B(abs_b[15]),
    .X(\v0/z4/z3/z3/temp [1]));
 sky130_fd_sc_hd__and2_0 \v0/z4/z3/z3/_3_  (.A(abs_a[9]),
    .B(abs_b[15]),
    .X(\v0/z4/z3/z3/temp [2]));
 sky130_fd_sc_hd__and2_0 \v0/z4/z3/z3/z1/_0_  (.A(\v0/z4/z3/z3/temp [1]),
    .B(\v0/z4/z3/z3/temp [0]),
    .X(\v0/z4/z3/z3/temp [3]));
 sky130_fd_sc_hd__xor2_1 \v0/z4/z3/z3/z1/_1_  (.A(\v0/z4/z3/z3/temp [1]),
    .B(\v0/z4/z3/z3/temp [0]),
    .X(\v0/z4/z3/q2 [1]));
 sky130_fd_sc_hd__and2_0 \v0/z4/z3/z3/z2/_0_  (.A(\v0/z4/z3/z3/temp [3]),
    .B(\v0/z4/z3/z3/temp [2]),
    .X(\v0/z4/z3/q2 [3]));
 sky130_fd_sc_hd__xor2_1 \v0/z4/z3/z3/z2/_1_  (.A(\v0/z4/z3/z3/temp [3]),
    .B(\v0/z4/z3/z3/temp [2]),
    .X(\v0/z4/z3/q2 [2]));
 sky130_fd_sc_hd__and2_0 \v0/z4/z3/z4/_0_  (.A(abs_b[14]),
    .B(abs_a[10]),
    .X(\v0/z4/z3/q3 [0]));
 sky130_fd_sc_hd__and2_0 \v0/z4/z3/z4/_1_  (.A(abs_b[14]),
    .B(abs_a[11]),
    .X(\v0/z4/z3/z4/temp [0]));
 sky130_fd_sc_hd__and2_0 \v0/z4/z3/z4/_2_  (.A(abs_a[10]),
    .B(abs_b[15]),
    .X(\v0/z4/z3/z4/temp [1]));
 sky130_fd_sc_hd__and2_0 \v0/z4/z3/z4/_3_  (.A(abs_a[11]),
    .B(abs_b[15]),
    .X(\v0/z4/z3/z4/temp [2]));
 sky130_fd_sc_hd__and2_0 \v0/z4/z3/z4/z1/_0_  (.A(\v0/z4/z3/z4/temp [1]),
    .B(\v0/z4/z3/z4/temp [0]),
    .X(\v0/z4/z3/z4/temp [3]));
 sky130_fd_sc_hd__xor2_1 \v0/z4/z3/z4/z1/_1_  (.A(\v0/z4/z3/z4/temp [1]),
    .B(\v0/z4/z3/z4/temp [0]),
    .X(\v0/z4/z3/q3 [1]));
 sky130_fd_sc_hd__and2_0 \v0/z4/z3/z4/z2/_0_  (.A(\v0/z4/z3/z4/temp [3]),
    .B(\v0/z4/z3/z4/temp [2]),
    .X(\v0/z4/z3/q3 [3]));
 sky130_fd_sc_hd__xor2_1 \v0/z4/z3/z4/z2/_1_  (.A(\v0/z4/z3/z4/temp [3]),
    .B(\v0/z4/z3/z4/temp [2]),
    .X(\v0/z4/z3/q3 [2]));
 sky130_fd_sc_hd__xnor2_1 \v0/z4/z3/z5/_07_  (.A(\v0/z4/z3/q0 [2]),
    .B(\v0/z4/z3/q1 [0]),
    .Y(\v0/z4/z3/z5/_00_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z4/z3/z5/_08_  (.A(\v0/z4/z3/_02_ ),
    .B(\v0/z4/z3/z5/_00_ ),
    .Y(\v0/z4/z3/q4 [0]));
 sky130_fd_sc_hd__maj3_1 \v0/z4/z3/z5/_09_  (.A(\v0/z4/z3/q0 [2]),
    .B(\v0/z4/z3/q1 [0]),
    .C(\v0/z4/z3/_02_ ),
    .X(\v0/z4/z3/z5/_01_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z4/z3/z5/_10_  (.A(\v0/z4/z3/q0 [3]),
    .B(\v0/z4/z3/q1 [1]),
    .Y(\v0/z4/z3/z5/_02_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z4/z3/z5/_11_  (.A(\v0/z4/z3/z5/_01_ ),
    .B(\v0/z4/z3/z5/_02_ ),
    .Y(\v0/z4/z3/q4 [1]));
 sky130_fd_sc_hd__maj3_1 \v0/z4/z3/z5/_12_  (.A(\v0/z4/z3/q0 [3]),
    .B(\v0/z4/z3/q1 [1]),
    .C(\v0/z4/z3/z5/_01_ ),
    .X(\v0/z4/z3/z5/_03_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z4/z3/z5/_13_  (.A(\v0/z4/z3/_00_ ),
    .B(\v0/z4/z3/q1 [2]),
    .Y(\v0/z4/z3/z5/_04_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z4/z3/z5/_14_  (.A(\v0/z4/z3/z5/_03_ ),
    .B(\v0/z4/z3/z5/_04_ ),
    .Y(\v0/z4/z3/q4 [2]));
 sky130_fd_sc_hd__maj3_1 \v0/z4/z3/z5/_15_  (.A(\v0/z4/z3/_00_ ),
    .B(\v0/z4/z3/q1 [2]),
    .C(\v0/z4/z3/z5/_03_ ),
    .X(\v0/z4/z3/z5/_05_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z4/z3/z5/_16_  (.A(\v0/z4/z3/_01_ ),
    .B(\v0/z4/z3/q1 [3]),
    .Y(\v0/z4/z3/z5/_06_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z4/z3/z5/_17_  (.A(\v0/z4/z3/z5/_05_ ),
    .B(\v0/z4/z3/z5/_06_ ),
    .Y(\v0/z4/z3/q4 [3]));
 sky130_fd_sc_hd__maj3_1 \v0/z4/z3/z5/_18_  (.A(\v0/z4/z3/_01_ ),
    .B(\v0/z4/z3/q1 [3]),
    .C(\v0/z4/z3/z5/_05_ ),
    .X(\v0/z4/z3/z5/Cout ));
 sky130_fd_sc_hd__xnor2_1 \v0/z4/z3/z6/_19_  (.A(\v0/z4/z3/_05_ ),
    .B(\v0/z4/z3/q2 [0]),
    .Y(\v0/z4/z3/z6/_00_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z4/z3/z6/_20_  (.A(\v0/z4/z3/_07_ ),
    .B(\v0/z4/z3/z6/_00_ ),
    .Y(\v0/z4/z3/q5 [0]));
 sky130_fd_sc_hd__maj3_1 \v0/z4/z3/z6/_21_  (.A(\v0/z4/z3/_05_ ),
    .B(\v0/z4/z3/q2 [0]),
    .C(\v0/z4/z3/_07_ ),
    .X(\v0/z4/z3/z6/_01_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z4/z3/z6/_22_  (.A(\v0/z4/z3/_06_ ),
    .B(\v0/z4/z3/q2 [1]),
    .Y(\v0/z4/z3/z6/_02_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z4/z3/z6/_23_  (.A(\v0/z4/z3/z6/_01_ ),
    .B(\v0/z4/z3/z6/_02_ ),
    .Y(\v0/z4/z3/q5 [1]));
 sky130_fd_sc_hd__maj3_1 \v0/z4/z3/z6/_24_  (.A(\v0/z4/z3/_06_ ),
    .B(\v0/z4/z3/q2 [1]),
    .C(\v0/z4/z3/z6/_01_ ),
    .X(\v0/z4/z3/z6/_03_ ));
 sky130_fd_sc_hd__lpflow_inputiso1p_1 \v0/z4/z3/z6/_25_  (.A(\v0/z4/z3/q3 [0]),
    .SLEEP(\v0/z4/z3/q2 [2]),
    .X(\v0/z4/z3/z6/_04_ ));
 sky130_fd_sc_hd__and2_0 \v0/z4/z3/z6/_26_  (.A(\v0/z4/z3/q3 [0]),
    .B(\v0/z4/z3/q2 [2]),
    .X(\v0/z4/z3/z6/_05_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z4/z3/z6/_27_  (.A(\v0/z4/z3/q3 [0]),
    .B(\v0/z4/z3/q2 [2]),
    .Y(\v0/z4/z3/z6/_06_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z4/z3/z6/_28_  (.A(\v0/z4/z3/z6/_04_ ),
    .B(\v0/z4/z3/z6/_06_ ),
    .Y(\v0/z4/z3/z6/_07_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z4/z3/z6/_29_  (.A(\v0/z4/z3/z6/_03_ ),
    .B(\v0/z4/z3/z6/_07_ ),
    .Y(\v0/z4/z3/q5 [2]));
 sky130_fd_sc_hd__nand2_1 \v0/z4/z3/z6/_30_  (.A(\v0/z4/z3/q3 [1]),
    .B(\v0/z4/z3/q2 [3]),
    .Y(\v0/z4/z3/z6/_08_ ));
 sky130_fd_sc_hd__xor2_1 \v0/z4/z3/z6/_31_  (.A(\v0/z4/z3/q3 [1]),
    .B(\v0/z4/z3/q2 [3]),
    .X(\v0/z4/z3/z6/_09_ ));
 sky130_fd_sc_hd__o21ai_0 \v0/z4/z3/z6/_32_  (.A1(\v0/z4/z3/z6/_03_ ),
    .A2(\v0/z4/z3/z6/_05_ ),
    .B1(\v0/z4/z3/z6/_04_ ),
    .Y(\v0/z4/z3/z6/_10_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z4/z3/z6/_33_  (.A(\v0/z4/z3/z6/_09_ ),
    .B(\v0/z4/z3/z6/_10_ ),
    .Y(\v0/z4/z3/q5 [3]));
 sky130_fd_sc_hd__nor2_1 \v0/z4/z3/z6/_34_  (.A(\v0/z4/z3/q3 [2]),
    .B(\v0/z4/z3/_03_ ),
    .Y(\v0/z4/z3/z6/_11_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z4/z3/z6/_35_  (.A(\v0/z4/z3/q3 [2]),
    .B(\v0/z4/z3/_03_ ),
    .Y(\v0/z4/z3/z6/_12_ ));
 sky130_fd_sc_hd__nand2b_1 \v0/z4/z3/z6/_36_  (.A_N(\v0/z4/z3/z6/_11_ ),
    .B(\v0/z4/z3/z6/_12_ ),
    .Y(\v0/z4/z3/z6/_13_ ));
 sky130_fd_sc_hd__o221ai_1 \v0/z4/z3/z6/_37_  (.A1(\v0/z4/z3/q3 [1]),
    .A2(\v0/z4/z3/q2 [3]),
    .B1(\v0/z4/z3/z6/_03_ ),
    .B2(\v0/z4/z3/z6/_05_ ),
    .C1(\v0/z4/z3/z6/_04_ ),
    .Y(\v0/z4/z3/z6/_14_ ));
 sky130_fd_sc_hd__a21oi_1 \v0/z4/z3/z6/_38_  (.A1(\v0/z4/z3/z6/_08_ ),
    .A2(\v0/z4/z3/z6/_14_ ),
    .B1(\v0/z4/z3/z6/_13_ ),
    .Y(\v0/z4/z3/z6/_15_ ));
 sky130_fd_sc_hd__and3_1 \v0/z4/z3/z6/_39_  (.A(\v0/z4/z3/z6/_08_ ),
    .B(\v0/z4/z3/z6/_13_ ),
    .C(\v0/z4/z3/z6/_14_ ),
    .X(\v0/z4/z3/z6/_16_ ));
 sky130_fd_sc_hd__nor2_1 \v0/z4/z3/z6/_40_  (.A(\v0/z4/z3/z6/_15_ ),
    .B(\v0/z4/z3/z6/_16_ ),
    .Y(\v0/z4/z3/q5 [4]));
 sky130_fd_sc_hd__xnor2_1 \v0/z4/z3/z6/_41_  (.A(\v0/z4/z3/q3 [3]),
    .B(\v0/z4/z3/_04_ ),
    .Y(\v0/z4/z3/z6/_17_ ));
 sky130_fd_sc_hd__a31oi_1 \v0/z4/z3/z6/_42_  (.A1(\v0/z4/z3/z6/_08_ ),
    .A2(\v0/z4/z3/z6/_12_ ),
    .A3(\v0/z4/z3/z6/_14_ ),
    .B1(\v0/z4/z3/z6/_11_ ),
    .Y(\v0/z4/z3/z6/_18_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z4/z3/z6/_43_  (.A(\v0/z4/z3/z6/_17_ ),
    .B(\v0/z4/z3/z6/_18_ ),
    .Y(\v0/z4/z3/q5 [5]));
 sky130_fd_sc_hd__maj3_1 \v0/z4/z3/z6/_44_  (.A(\v0/z4/z3/q3 [3]),
    .B(\v0/z4/z3/_04_ ),
    .C(\v0/z4/z3/z6/_18_ ),
    .X(\v0/z4/z3/z6/Cout ));
 sky130_fd_sc_hd__xnor2_1 \v0/z4/z3/z7/_19_  (.A(\v0/z4/z3/q5 [0]),
    .B(\v0/z4/z3/q4 [0]),
    .Y(\v0/z4/z3/z7/_00_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z4/z3/z7/_20_  (.A(\v0/z4/z3/_10_ ),
    .B(\v0/z4/z3/z7/_00_ ),
    .Y(\v0/z4/q2 [2]));
 sky130_fd_sc_hd__maj3_1 \v0/z4/z3/z7/_21_  (.A(\v0/z4/z3/q5 [0]),
    .B(\v0/z4/z3/q4 [0]),
    .C(\v0/z4/z3/_10_ ),
    .X(\v0/z4/z3/z7/_01_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z4/z3/z7/_22_  (.A(\v0/z4/z3/q5 [1]),
    .B(\v0/z4/z3/q4 [1]),
    .Y(\v0/z4/z3/z7/_02_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z4/z3/z7/_23_  (.A(\v0/z4/z3/z7/_01_ ),
    .B(\v0/z4/z3/z7/_02_ ),
    .Y(\v0/z4/q2 [3]));
 sky130_fd_sc_hd__maj3_1 \v0/z4/z3/z7/_24_  (.A(\v0/z4/z3/q5 [1]),
    .B(\v0/z4/z3/q4 [1]),
    .C(\v0/z4/z3/z7/_01_ ),
    .X(\v0/z4/z3/z7/_03_ ));
 sky130_fd_sc_hd__lpflow_inputiso1p_1 \v0/z4/z3/z7/_25_  (.A(\v0/z4/z3/q5 [2]),
    .SLEEP(\v0/z4/z3/q4 [2]),
    .X(\v0/z4/z3/z7/_04_ ));
 sky130_fd_sc_hd__and2_0 \v0/z4/z3/z7/_26_  (.A(\v0/z4/z3/q5 [2]),
    .B(\v0/z4/z3/q4 [2]),
    .X(\v0/z4/z3/z7/_05_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z4/z3/z7/_27_  (.A(\v0/z4/z3/q5 [2]),
    .B(\v0/z4/z3/q4 [2]),
    .Y(\v0/z4/z3/z7/_06_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z4/z3/z7/_28_  (.A(\v0/z4/z3/z7/_04_ ),
    .B(\v0/z4/z3/z7/_06_ ),
    .Y(\v0/z4/z3/z7/_07_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z4/z3/z7/_29_  (.A(\v0/z4/z3/z7/_03_ ),
    .B(\v0/z4/z3/z7/_07_ ),
    .Y(\v0/z4/q2 [4]));
 sky130_fd_sc_hd__nand2_1 \v0/z4/z3/z7/_30_  (.A(\v0/z4/z3/q5 [3]),
    .B(\v0/z4/z3/q4 [3]),
    .Y(\v0/z4/z3/z7/_08_ ));
 sky130_fd_sc_hd__xor2_1 \v0/z4/z3/z7/_31_  (.A(\v0/z4/z3/q5 [3]),
    .B(\v0/z4/z3/q4 [3]),
    .X(\v0/z4/z3/z7/_09_ ));
 sky130_fd_sc_hd__o21ai_0 \v0/z4/z3/z7/_32_  (.A1(\v0/z4/z3/z7/_03_ ),
    .A2(\v0/z4/z3/z7/_05_ ),
    .B1(\v0/z4/z3/z7/_04_ ),
    .Y(\v0/z4/z3/z7/_10_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z4/z3/z7/_33_  (.A(\v0/z4/z3/z7/_09_ ),
    .B(\v0/z4/z3/z7/_10_ ),
    .Y(\v0/z4/q2 [5]));
 sky130_fd_sc_hd__nor2_1 \v0/z4/z3/z7/_34_  (.A(\v0/z4/z3/q5 [4]),
    .B(\v0/z4/z3/_08_ ),
    .Y(\v0/z4/z3/z7/_11_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z4/z3/z7/_35_  (.A(\v0/z4/z3/q5 [4]),
    .B(\v0/z4/z3/_08_ ),
    .Y(\v0/z4/z3/z7/_12_ ));
 sky130_fd_sc_hd__nand2b_1 \v0/z4/z3/z7/_36_  (.A_N(\v0/z4/z3/z7/_11_ ),
    .B(\v0/z4/z3/z7/_12_ ),
    .Y(\v0/z4/z3/z7/_13_ ));
 sky130_fd_sc_hd__o221ai_1 \v0/z4/z3/z7/_37_  (.A1(\v0/z4/z3/q5 [3]),
    .A2(\v0/z4/z3/q4 [3]),
    .B1(\v0/z4/z3/z7/_03_ ),
    .B2(\v0/z4/z3/z7/_05_ ),
    .C1(\v0/z4/z3/z7/_04_ ),
    .Y(\v0/z4/z3/z7/_14_ ));
 sky130_fd_sc_hd__a21oi_1 \v0/z4/z3/z7/_38_  (.A1(\v0/z4/z3/z7/_08_ ),
    .A2(\v0/z4/z3/z7/_14_ ),
    .B1(\v0/z4/z3/z7/_13_ ),
    .Y(\v0/z4/z3/z7/_15_ ));
 sky130_fd_sc_hd__and3_1 \v0/z4/z3/z7/_39_  (.A(\v0/z4/z3/z7/_08_ ),
    .B(\v0/z4/z3/z7/_13_ ),
    .C(\v0/z4/z3/z7/_14_ ),
    .X(\v0/z4/z3/z7/_16_ ));
 sky130_fd_sc_hd__nor2_1 \v0/z4/z3/z7/_40_  (.A(\v0/z4/z3/z7/_15_ ),
    .B(\v0/z4/z3/z7/_16_ ),
    .Y(\v0/z4/q2 [6]));
 sky130_fd_sc_hd__xnor2_1 \v0/z4/z3/z7/_41_  (.A(\v0/z4/z3/q5 [5]),
    .B(\v0/z4/z3/_09_ ),
    .Y(\v0/z4/z3/z7/_17_ ));
 sky130_fd_sc_hd__a31oi_1 \v0/z4/z3/z7/_42_  (.A1(\v0/z4/z3/z7/_08_ ),
    .A2(\v0/z4/z3/z7/_12_ ),
    .A3(\v0/z4/z3/z7/_14_ ),
    .B1(\v0/z4/z3/z7/_11_ ),
    .Y(\v0/z4/z3/z7/_18_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z4/z3/z7/_43_  (.A(\v0/z4/z3/z7/_17_ ),
    .B(\v0/z4/z3/z7/_18_ ),
    .Y(\v0/z4/q2 [7]));
 sky130_fd_sc_hd__maj3_1 \v0/z4/z3/z7/_44_  (.A(\v0/z4/z3/q5 [5]),
    .B(\v0/z4/z3/_09_ ),
    .C(\v0/z4/z3/z7/_18_ ),
    .X(\v0/z4/z3/z7/Cout ));
 sky130_fd_sc_hd__conb_1 \v0/z4/z4/_11_  (.LO(\v0/z4/z4/_00_ ));
 sky130_fd_sc_hd__conb_1 \v0/z4/z4/_12_  (.LO(\v0/z4/z4/_01_ ));
 sky130_fd_sc_hd__conb_1 \v0/z4/z4/_13_  (.LO(\v0/z4/z4/_02_ ));
 sky130_fd_sc_hd__conb_1 \v0/z4/z4/_14_  (.LO(\v0/z4/z4/_03_ ));
 sky130_fd_sc_hd__conb_1 \v0/z4/z4/_15_  (.LO(\v0/z4/z4/_04_ ));
 sky130_fd_sc_hd__conb_1 \v0/z4/z4/_16_  (.LO(\v0/z4/z4/_05_ ));
 sky130_fd_sc_hd__conb_1 \v0/z4/z4/_17_  (.LO(\v0/z4/z4/_06_ ));
 sky130_fd_sc_hd__conb_1 \v0/z4/z4/_18_  (.LO(\v0/z4/z4/_07_ ));
 sky130_fd_sc_hd__conb_1 \v0/z4/z4/_19_  (.LO(\v0/z4/z4/_08_ ));
 sky130_fd_sc_hd__conb_1 \v0/z4/z4/_20_  (.LO(\v0/z4/z4/_09_ ));
 sky130_fd_sc_hd__conb_1 \v0/z4/z4/_21_  (.LO(\v0/z4/z4/_10_ ));
 sky130_fd_sc_hd__and2_0 \v0/z4/z4/z1/_0_  (.A(abs_b[12]),
    .B(abs_a[12]),
    .X(\v0/z4/q3 [0]));
 sky130_fd_sc_hd__and2_0 \v0/z4/z4/z1/_1_  (.A(abs_b[12]),
    .B(abs_a[13]),
    .X(\v0/z4/z4/z1/temp [0]));
 sky130_fd_sc_hd__and2_0 \v0/z4/z4/z1/_2_  (.A(abs_a[12]),
    .B(abs_b[13]),
    .X(\v0/z4/z4/z1/temp [1]));
 sky130_fd_sc_hd__and2_0 \v0/z4/z4/z1/_3_  (.A(abs_a[13]),
    .B(abs_b[13]),
    .X(\v0/z4/z4/z1/temp [2]));
 sky130_fd_sc_hd__and2_0 \v0/z4/z4/z1/z1/_0_  (.A(\v0/z4/z4/z1/temp [1]),
    .B(\v0/z4/z4/z1/temp [0]),
    .X(\v0/z4/z4/z1/temp [3]));
 sky130_fd_sc_hd__xor2_1 \v0/z4/z4/z1/z1/_1_  (.A(\v0/z4/z4/z1/temp [1]),
    .B(\v0/z4/z4/z1/temp [0]),
    .X(\v0/z4/q3 [1]));
 sky130_fd_sc_hd__and2_0 \v0/z4/z4/z1/z2/_0_  (.A(\v0/z4/z4/z1/temp [3]),
    .B(\v0/z4/z4/z1/temp [2]),
    .X(\v0/z4/z4/q0 [3]));
 sky130_fd_sc_hd__xor2_1 \v0/z4/z4/z1/z2/_1_  (.A(\v0/z4/z4/z1/temp [3]),
    .B(\v0/z4/z4/z1/temp [2]),
    .X(\v0/z4/z4/q0 [2]));
 sky130_fd_sc_hd__and2_0 \v0/z4/z4/z2/_0_  (.A(abs_b[12]),
    .B(abs_a[14]),
    .X(\v0/z4/z4/q1 [0]));
 sky130_fd_sc_hd__and2_0 \v0/z4/z4/z2/_1_  (.A(abs_b[12]),
    .B(abs_a[15]),
    .X(\v0/z4/z4/z2/temp [0]));
 sky130_fd_sc_hd__and2_0 \v0/z4/z4/z2/_2_  (.A(abs_a[14]),
    .B(abs_b[13]),
    .X(\v0/z4/z4/z2/temp [1]));
 sky130_fd_sc_hd__and2_0 \v0/z4/z4/z2/_3_  (.A(abs_a[15]),
    .B(abs_b[13]),
    .X(\v0/z4/z4/z2/temp [2]));
 sky130_fd_sc_hd__and2_0 \v0/z4/z4/z2/z1/_0_  (.A(\v0/z4/z4/z2/temp [1]),
    .B(\v0/z4/z4/z2/temp [0]),
    .X(\v0/z4/z4/z2/temp [3]));
 sky130_fd_sc_hd__xor2_1 \v0/z4/z4/z2/z1/_1_  (.A(\v0/z4/z4/z2/temp [1]),
    .B(\v0/z4/z4/z2/temp [0]),
    .X(\v0/z4/z4/q1 [1]));
 sky130_fd_sc_hd__and2_0 \v0/z4/z4/z2/z2/_0_  (.A(\v0/z4/z4/z2/temp [3]),
    .B(\v0/z4/z4/z2/temp [2]),
    .X(\v0/z4/z4/q1 [3]));
 sky130_fd_sc_hd__xor2_1 \v0/z4/z4/z2/z2/_1_  (.A(\v0/z4/z4/z2/temp [3]),
    .B(\v0/z4/z4/z2/temp [2]),
    .X(\v0/z4/z4/q1 [2]));
 sky130_fd_sc_hd__and2_0 \v0/z4/z4/z3/_0_  (.A(abs_b[14]),
    .B(abs_a[12]),
    .X(\v0/z4/z4/q2 [0]));
 sky130_fd_sc_hd__and2_0 \v0/z4/z4/z3/_1_  (.A(abs_b[14]),
    .B(abs_a[13]),
    .X(\v0/z4/z4/z3/temp [0]));
 sky130_fd_sc_hd__and2_0 \v0/z4/z4/z3/_2_  (.A(abs_a[12]),
    .B(abs_b[15]),
    .X(\v0/z4/z4/z3/temp [1]));
 sky130_fd_sc_hd__and2_0 \v0/z4/z4/z3/_3_  (.A(abs_a[13]),
    .B(abs_b[15]),
    .X(\v0/z4/z4/z3/temp [2]));
 sky130_fd_sc_hd__and2_0 \v0/z4/z4/z3/z1/_0_  (.A(\v0/z4/z4/z3/temp [1]),
    .B(\v0/z4/z4/z3/temp [0]),
    .X(\v0/z4/z4/z3/temp [3]));
 sky130_fd_sc_hd__xor2_1 \v0/z4/z4/z3/z1/_1_  (.A(\v0/z4/z4/z3/temp [1]),
    .B(\v0/z4/z4/z3/temp [0]),
    .X(\v0/z4/z4/q2 [1]));
 sky130_fd_sc_hd__and2_0 \v0/z4/z4/z3/z2/_0_  (.A(\v0/z4/z4/z3/temp [3]),
    .B(\v0/z4/z4/z3/temp [2]),
    .X(\v0/z4/z4/q2 [3]));
 sky130_fd_sc_hd__xor2_1 \v0/z4/z4/z3/z2/_1_  (.A(\v0/z4/z4/z3/temp [3]),
    .B(\v0/z4/z4/z3/temp [2]),
    .X(\v0/z4/z4/q2 [2]));
 sky130_fd_sc_hd__and2_0 \v0/z4/z4/z4/_0_  (.A(abs_b[14]),
    .B(abs_a[14]),
    .X(\v0/z4/z4/q3 [0]));
 sky130_fd_sc_hd__and2_0 \v0/z4/z4/z4/_1_  (.A(abs_b[14]),
    .B(abs_a[15]),
    .X(\v0/z4/z4/z4/temp [0]));
 sky130_fd_sc_hd__and2_0 \v0/z4/z4/z4/_2_  (.A(abs_a[14]),
    .B(abs_b[15]),
    .X(\v0/z4/z4/z4/temp [1]));
 sky130_fd_sc_hd__and2_0 \v0/z4/z4/z4/_3_  (.A(abs_a[15]),
    .B(abs_b[15]),
    .X(\v0/z4/z4/z4/temp [2]));
 sky130_fd_sc_hd__and2_0 \v0/z4/z4/z4/z1/_0_  (.A(\v0/z4/z4/z4/temp [1]),
    .B(\v0/z4/z4/z4/temp [0]),
    .X(\v0/z4/z4/z4/temp [3]));
 sky130_fd_sc_hd__xor2_1 \v0/z4/z4/z4/z1/_1_  (.A(\v0/z4/z4/z4/temp [1]),
    .B(\v0/z4/z4/z4/temp [0]),
    .X(\v0/z4/z4/q3 [1]));
 sky130_fd_sc_hd__and2_0 \v0/z4/z4/z4/z2/_0_  (.A(\v0/z4/z4/z4/temp [3]),
    .B(\v0/z4/z4/z4/temp [2]),
    .X(\v0/z4/z4/q3 [3]));
 sky130_fd_sc_hd__xor2_1 \v0/z4/z4/z4/z2/_1_  (.A(\v0/z4/z4/z4/temp [3]),
    .B(\v0/z4/z4/z4/temp [2]),
    .X(\v0/z4/z4/q3 [2]));
 sky130_fd_sc_hd__xnor2_1 \v0/z4/z4/z5/_07_  (.A(\v0/z4/z4/q0 [2]),
    .B(\v0/z4/z4/q1 [0]),
    .Y(\v0/z4/z4/z5/_00_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z4/z4/z5/_08_  (.A(\v0/z4/z4/_02_ ),
    .B(\v0/z4/z4/z5/_00_ ),
    .Y(\v0/z4/z4/q4 [0]));
 sky130_fd_sc_hd__maj3_1 \v0/z4/z4/z5/_09_  (.A(\v0/z4/z4/q0 [2]),
    .B(\v0/z4/z4/q1 [0]),
    .C(\v0/z4/z4/_02_ ),
    .X(\v0/z4/z4/z5/_01_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z4/z4/z5/_10_  (.A(\v0/z4/z4/q0 [3]),
    .B(\v0/z4/z4/q1 [1]),
    .Y(\v0/z4/z4/z5/_02_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z4/z4/z5/_11_  (.A(\v0/z4/z4/z5/_01_ ),
    .B(\v0/z4/z4/z5/_02_ ),
    .Y(\v0/z4/z4/q4 [1]));
 sky130_fd_sc_hd__maj3_1 \v0/z4/z4/z5/_12_  (.A(\v0/z4/z4/q0 [3]),
    .B(\v0/z4/z4/q1 [1]),
    .C(\v0/z4/z4/z5/_01_ ),
    .X(\v0/z4/z4/z5/_03_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z4/z4/z5/_13_  (.A(\v0/z4/z4/_00_ ),
    .B(\v0/z4/z4/q1 [2]),
    .Y(\v0/z4/z4/z5/_04_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z4/z4/z5/_14_  (.A(\v0/z4/z4/z5/_03_ ),
    .B(\v0/z4/z4/z5/_04_ ),
    .Y(\v0/z4/z4/q4 [2]));
 sky130_fd_sc_hd__maj3_1 \v0/z4/z4/z5/_15_  (.A(\v0/z4/z4/_00_ ),
    .B(\v0/z4/z4/q1 [2]),
    .C(\v0/z4/z4/z5/_03_ ),
    .X(\v0/z4/z4/z5/_05_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z4/z4/z5/_16_  (.A(\v0/z4/z4/_01_ ),
    .B(\v0/z4/z4/q1 [3]),
    .Y(\v0/z4/z4/z5/_06_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z4/z4/z5/_17_  (.A(\v0/z4/z4/z5/_05_ ),
    .B(\v0/z4/z4/z5/_06_ ),
    .Y(\v0/z4/z4/q4 [3]));
 sky130_fd_sc_hd__maj3_1 \v0/z4/z4/z5/_18_  (.A(\v0/z4/z4/_01_ ),
    .B(\v0/z4/z4/q1 [3]),
    .C(\v0/z4/z4/z5/_05_ ),
    .X(\v0/z4/z4/z5/Cout ));
 sky130_fd_sc_hd__xnor2_1 \v0/z4/z4/z6/_19_  (.A(\v0/z4/z4/_05_ ),
    .B(\v0/z4/z4/q2 [0]),
    .Y(\v0/z4/z4/z6/_00_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z4/z4/z6/_20_  (.A(\v0/z4/z4/_07_ ),
    .B(\v0/z4/z4/z6/_00_ ),
    .Y(\v0/z4/z4/q5 [0]));
 sky130_fd_sc_hd__maj3_1 \v0/z4/z4/z6/_21_  (.A(\v0/z4/z4/_05_ ),
    .B(\v0/z4/z4/q2 [0]),
    .C(\v0/z4/z4/_07_ ),
    .X(\v0/z4/z4/z6/_01_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z4/z4/z6/_22_  (.A(\v0/z4/z4/_06_ ),
    .B(\v0/z4/z4/q2 [1]),
    .Y(\v0/z4/z4/z6/_02_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z4/z4/z6/_23_  (.A(\v0/z4/z4/z6/_01_ ),
    .B(\v0/z4/z4/z6/_02_ ),
    .Y(\v0/z4/z4/q5 [1]));
 sky130_fd_sc_hd__maj3_1 \v0/z4/z4/z6/_24_  (.A(\v0/z4/z4/_06_ ),
    .B(\v0/z4/z4/q2 [1]),
    .C(\v0/z4/z4/z6/_01_ ),
    .X(\v0/z4/z4/z6/_03_ ));
 sky130_fd_sc_hd__lpflow_inputiso1p_1 \v0/z4/z4/z6/_25_  (.A(\v0/z4/z4/q3 [0]),
    .SLEEP(\v0/z4/z4/q2 [2]),
    .X(\v0/z4/z4/z6/_04_ ));
 sky130_fd_sc_hd__and2_0 \v0/z4/z4/z6/_26_  (.A(\v0/z4/z4/q3 [0]),
    .B(\v0/z4/z4/q2 [2]),
    .X(\v0/z4/z4/z6/_05_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z4/z4/z6/_27_  (.A(\v0/z4/z4/q3 [0]),
    .B(\v0/z4/z4/q2 [2]),
    .Y(\v0/z4/z4/z6/_06_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z4/z4/z6/_28_  (.A(\v0/z4/z4/z6/_04_ ),
    .B(\v0/z4/z4/z6/_06_ ),
    .Y(\v0/z4/z4/z6/_07_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z4/z4/z6/_29_  (.A(\v0/z4/z4/z6/_03_ ),
    .B(\v0/z4/z4/z6/_07_ ),
    .Y(\v0/z4/z4/q5 [2]));
 sky130_fd_sc_hd__nand2_1 \v0/z4/z4/z6/_30_  (.A(\v0/z4/z4/q3 [1]),
    .B(\v0/z4/z4/q2 [3]),
    .Y(\v0/z4/z4/z6/_08_ ));
 sky130_fd_sc_hd__xor2_1 \v0/z4/z4/z6/_31_  (.A(\v0/z4/z4/q3 [1]),
    .B(\v0/z4/z4/q2 [3]),
    .X(\v0/z4/z4/z6/_09_ ));
 sky130_fd_sc_hd__o21ai_0 \v0/z4/z4/z6/_32_  (.A1(\v0/z4/z4/z6/_03_ ),
    .A2(\v0/z4/z4/z6/_05_ ),
    .B1(\v0/z4/z4/z6/_04_ ),
    .Y(\v0/z4/z4/z6/_10_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z4/z4/z6/_33_  (.A(\v0/z4/z4/z6/_09_ ),
    .B(\v0/z4/z4/z6/_10_ ),
    .Y(\v0/z4/z4/q5 [3]));
 sky130_fd_sc_hd__nor2_1 \v0/z4/z4/z6/_34_  (.A(\v0/z4/z4/q3 [2]),
    .B(\v0/z4/z4/_03_ ),
    .Y(\v0/z4/z4/z6/_11_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z4/z4/z6/_35_  (.A(\v0/z4/z4/q3 [2]),
    .B(\v0/z4/z4/_03_ ),
    .Y(\v0/z4/z4/z6/_12_ ));
 sky130_fd_sc_hd__nand2b_1 \v0/z4/z4/z6/_36_  (.A_N(\v0/z4/z4/z6/_11_ ),
    .B(\v0/z4/z4/z6/_12_ ),
    .Y(\v0/z4/z4/z6/_13_ ));
 sky130_fd_sc_hd__o221ai_1 \v0/z4/z4/z6/_37_  (.A1(\v0/z4/z4/q3 [1]),
    .A2(\v0/z4/z4/q2 [3]),
    .B1(\v0/z4/z4/z6/_03_ ),
    .B2(\v0/z4/z4/z6/_05_ ),
    .C1(\v0/z4/z4/z6/_04_ ),
    .Y(\v0/z4/z4/z6/_14_ ));
 sky130_fd_sc_hd__a21oi_1 \v0/z4/z4/z6/_38_  (.A1(\v0/z4/z4/z6/_08_ ),
    .A2(\v0/z4/z4/z6/_14_ ),
    .B1(\v0/z4/z4/z6/_13_ ),
    .Y(\v0/z4/z4/z6/_15_ ));
 sky130_fd_sc_hd__and3_1 \v0/z4/z4/z6/_39_  (.A(\v0/z4/z4/z6/_08_ ),
    .B(\v0/z4/z4/z6/_13_ ),
    .C(\v0/z4/z4/z6/_14_ ),
    .X(\v0/z4/z4/z6/_16_ ));
 sky130_fd_sc_hd__nor2_1 \v0/z4/z4/z6/_40_  (.A(\v0/z4/z4/z6/_15_ ),
    .B(\v0/z4/z4/z6/_16_ ),
    .Y(\v0/z4/z4/q5 [4]));
 sky130_fd_sc_hd__xnor2_1 \v0/z4/z4/z6/_41_  (.A(\v0/z4/z4/q3 [3]),
    .B(\v0/z4/z4/_04_ ),
    .Y(\v0/z4/z4/z6/_17_ ));
 sky130_fd_sc_hd__a31oi_1 \v0/z4/z4/z6/_42_  (.A1(\v0/z4/z4/z6/_08_ ),
    .A2(\v0/z4/z4/z6/_12_ ),
    .A3(\v0/z4/z4/z6/_14_ ),
    .B1(\v0/z4/z4/z6/_11_ ),
    .Y(\v0/z4/z4/z6/_18_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z4/z4/z6/_43_  (.A(\v0/z4/z4/z6/_17_ ),
    .B(\v0/z4/z4/z6/_18_ ),
    .Y(\v0/z4/z4/q5 [5]));
 sky130_fd_sc_hd__maj3_1 \v0/z4/z4/z6/_44_  (.A(\v0/z4/z4/q3 [3]),
    .B(\v0/z4/z4/_04_ ),
    .C(\v0/z4/z4/z6/_18_ ),
    .X(\v0/z4/z4/z6/Cout ));
 sky130_fd_sc_hd__xnor2_1 \v0/z4/z4/z7/_19_  (.A(\v0/z4/z4/q5 [0]),
    .B(\v0/z4/z4/q4 [0]),
    .Y(\v0/z4/z4/z7/_00_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z4/z4/z7/_20_  (.A(\v0/z4/z4/_10_ ),
    .B(\v0/z4/z4/z7/_00_ ),
    .Y(\v0/z4/q3 [2]));
 sky130_fd_sc_hd__maj3_1 \v0/z4/z4/z7/_21_  (.A(\v0/z4/z4/q5 [0]),
    .B(\v0/z4/z4/q4 [0]),
    .C(\v0/z4/z4/_10_ ),
    .X(\v0/z4/z4/z7/_01_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z4/z4/z7/_22_  (.A(\v0/z4/z4/q5 [1]),
    .B(\v0/z4/z4/q4 [1]),
    .Y(\v0/z4/z4/z7/_02_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z4/z4/z7/_23_  (.A(\v0/z4/z4/z7/_01_ ),
    .B(\v0/z4/z4/z7/_02_ ),
    .Y(\v0/z4/q3 [3]));
 sky130_fd_sc_hd__maj3_1 \v0/z4/z4/z7/_24_  (.A(\v0/z4/z4/q5 [1]),
    .B(\v0/z4/z4/q4 [1]),
    .C(\v0/z4/z4/z7/_01_ ),
    .X(\v0/z4/z4/z7/_03_ ));
 sky130_fd_sc_hd__lpflow_inputiso1p_1 \v0/z4/z4/z7/_25_  (.A(\v0/z4/z4/q5 [2]),
    .SLEEP(\v0/z4/z4/q4 [2]),
    .X(\v0/z4/z4/z7/_04_ ));
 sky130_fd_sc_hd__and2_0 \v0/z4/z4/z7/_26_  (.A(\v0/z4/z4/q5 [2]),
    .B(\v0/z4/z4/q4 [2]),
    .X(\v0/z4/z4/z7/_05_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z4/z4/z7/_27_  (.A(\v0/z4/z4/q5 [2]),
    .B(\v0/z4/z4/q4 [2]),
    .Y(\v0/z4/z4/z7/_06_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z4/z4/z7/_28_  (.A(\v0/z4/z4/z7/_04_ ),
    .B(\v0/z4/z4/z7/_06_ ),
    .Y(\v0/z4/z4/z7/_07_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z4/z4/z7/_29_  (.A(\v0/z4/z4/z7/_03_ ),
    .B(\v0/z4/z4/z7/_07_ ),
    .Y(\v0/z4/q3 [4]));
 sky130_fd_sc_hd__nand2_1 \v0/z4/z4/z7/_30_  (.A(\v0/z4/z4/q5 [3]),
    .B(\v0/z4/z4/q4 [3]),
    .Y(\v0/z4/z4/z7/_08_ ));
 sky130_fd_sc_hd__xor2_1 \v0/z4/z4/z7/_31_  (.A(\v0/z4/z4/q5 [3]),
    .B(\v0/z4/z4/q4 [3]),
    .X(\v0/z4/z4/z7/_09_ ));
 sky130_fd_sc_hd__o21ai_0 \v0/z4/z4/z7/_32_  (.A1(\v0/z4/z4/z7/_03_ ),
    .A2(\v0/z4/z4/z7/_05_ ),
    .B1(\v0/z4/z4/z7/_04_ ),
    .Y(\v0/z4/z4/z7/_10_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z4/z4/z7/_33_  (.A(\v0/z4/z4/z7/_09_ ),
    .B(\v0/z4/z4/z7/_10_ ),
    .Y(\v0/z4/q3 [5]));
 sky130_fd_sc_hd__nor2_1 \v0/z4/z4/z7/_34_  (.A(\v0/z4/z4/q5 [4]),
    .B(\v0/z4/z4/_08_ ),
    .Y(\v0/z4/z4/z7/_11_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z4/z4/z7/_35_  (.A(\v0/z4/z4/q5 [4]),
    .B(\v0/z4/z4/_08_ ),
    .Y(\v0/z4/z4/z7/_12_ ));
 sky130_fd_sc_hd__nand2b_1 \v0/z4/z4/z7/_36_  (.A_N(\v0/z4/z4/z7/_11_ ),
    .B(\v0/z4/z4/z7/_12_ ),
    .Y(\v0/z4/z4/z7/_13_ ));
 sky130_fd_sc_hd__o221ai_1 \v0/z4/z4/z7/_37_  (.A1(\v0/z4/z4/q5 [3]),
    .A2(\v0/z4/z4/q4 [3]),
    .B1(\v0/z4/z4/z7/_03_ ),
    .B2(\v0/z4/z4/z7/_05_ ),
    .C1(\v0/z4/z4/z7/_04_ ),
    .Y(\v0/z4/z4/z7/_14_ ));
 sky130_fd_sc_hd__a21oi_1 \v0/z4/z4/z7/_38_  (.A1(\v0/z4/z4/z7/_08_ ),
    .A2(\v0/z4/z4/z7/_14_ ),
    .B1(\v0/z4/z4/z7/_13_ ),
    .Y(\v0/z4/z4/z7/_15_ ));
 sky130_fd_sc_hd__and3_1 \v0/z4/z4/z7/_39_  (.A(\v0/z4/z4/z7/_08_ ),
    .B(\v0/z4/z4/z7/_13_ ),
    .C(\v0/z4/z4/z7/_14_ ),
    .X(\v0/z4/z4/z7/_16_ ));
 sky130_fd_sc_hd__nor2_1 \v0/z4/z4/z7/_40_  (.A(\v0/z4/z4/z7/_15_ ),
    .B(\v0/z4/z4/z7/_16_ ),
    .Y(\v0/z4/q3 [6]));
 sky130_fd_sc_hd__xnor2_1 \v0/z4/z4/z7/_41_  (.A(\v0/z4/z4/q5 [5]),
    .B(\v0/z4/z4/_09_ ),
    .Y(\v0/z4/z4/z7/_17_ ));
 sky130_fd_sc_hd__a31oi_1 \v0/z4/z4/z7/_42_  (.A1(\v0/z4/z4/z7/_08_ ),
    .A2(\v0/z4/z4/z7/_12_ ),
    .A3(\v0/z4/z4/z7/_14_ ),
    .B1(\v0/z4/z4/z7/_11_ ),
    .Y(\v0/z4/z4/z7/_18_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z4/z4/z7/_43_  (.A(\v0/z4/z4/z7/_17_ ),
    .B(\v0/z4/z4/z7/_18_ ),
    .Y(\v0/z4/q3 [7]));
 sky130_fd_sc_hd__maj3_1 \v0/z4/z4/z7/_44_  (.A(\v0/z4/z4/q5 [5]),
    .B(\v0/z4/z4/_09_ ),
    .C(\v0/z4/z4/z7/_18_ ),
    .X(\v0/z4/z4/z7/Cout ));
 sky130_fd_sc_hd__xnor2_1 \v0/z4/z5/_27_  (.A(\v0/z4/q0 [4]),
    .B(\v0/z4/q1 [0]),
    .Y(\v0/z4/z5/_00_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z4/z5/_28_  (.A(\v0/z4/_04_ ),
    .B(\v0/z4/z5/_00_ ),
    .Y(\v0/z4/q4 [0]));
 sky130_fd_sc_hd__maj3_1 \v0/z4/z5/_29_  (.A(\v0/z4/q0 [4]),
    .B(\v0/z4/q1 [0]),
    .C(\v0/z4/_04_ ),
    .X(\v0/z4/z5/_01_ ));
 sky130_fd_sc_hd__lpflow_inputiso1p_1 \v0/z4/z5/_30_  (.A(\v0/z4/q0 [5]),
    .SLEEP(\v0/z4/q1 [1]),
    .X(\v0/z4/z5/_02_ ));
 sky130_fd_sc_hd__and2_0 \v0/z4/z5/_31_  (.A(\v0/z4/q0 [5]),
    .B(\v0/z4/q1 [1]),
    .X(\v0/z4/z5/_03_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z4/z5/_32_  (.A(\v0/z4/q0 [5]),
    .B(\v0/z4/q1 [1]),
    .Y(\v0/z4/z5/_04_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z4/z5/_33_  (.A(\v0/z4/z5/_02_ ),
    .B(\v0/z4/z5/_04_ ),
    .Y(\v0/z4/z5/_05_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z4/z5/_34_  (.A(\v0/z4/z5/_01_ ),
    .B(\v0/z4/z5/_05_ ),
    .Y(\v0/z4/q4 [1]));
 sky130_fd_sc_hd__nand2_1 \v0/z4/z5/_35_  (.A(\v0/z4/q0 [6]),
    .B(\v0/z4/q1 [2]),
    .Y(\v0/z4/z5/_06_ ));
 sky130_fd_sc_hd__xor2_1 \v0/z4/z5/_36_  (.A(\v0/z4/q0 [6]),
    .B(\v0/z4/q1 [2]),
    .X(\v0/z4/z5/_07_ ));
 sky130_fd_sc_hd__o21ai_0 \v0/z4/z5/_37_  (.A1(\v0/z4/z5/_01_ ),
    .A2(\v0/z4/z5/_03_ ),
    .B1(\v0/z4/z5/_02_ ),
    .Y(\v0/z4/z5/_08_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z4/z5/_38_  (.A(\v0/z4/z5/_07_ ),
    .B(\v0/z4/z5/_08_ ),
    .Y(\v0/z4/q4 [2]));
 sky130_fd_sc_hd__nor2_1 \v0/z4/z5/_39_  (.A(\v0/z4/q0 [7]),
    .B(\v0/z4/q1 [3]),
    .Y(\v0/z4/z5/_09_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z4/z5/_40_  (.A(\v0/z4/q0 [7]),
    .B(\v0/z4/q1 [3]),
    .Y(\v0/z4/z5/_10_ ));
 sky130_fd_sc_hd__nor2b_1 \v0/z4/z5/_41_  (.A(\v0/z4/z5/_09_ ),
    .B_N(\v0/z4/z5/_10_ ),
    .Y(\v0/z4/z5/_11_ ));
 sky130_fd_sc_hd__o221ai_1 \v0/z4/z5/_42_  (.A1(\v0/z4/q0 [6]),
    .A2(\v0/z4/q1 [2]),
    .B1(\v0/z4/z5/_01_ ),
    .B2(\v0/z4/z5/_03_ ),
    .C1(\v0/z4/z5/_02_ ),
    .Y(\v0/z4/z5/_12_ ));
 sky130_fd_sc_hd__and2_0 \v0/z4/z5/_43_  (.A(\v0/z4/z5/_06_ ),
    .B(\v0/z4/z5/_12_ ),
    .X(\v0/z4/z5/_13_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z4/z5/_44_  (.A(\v0/z4/z5/_11_ ),
    .B(\v0/z4/z5/_13_ ),
    .Y(\v0/z4/q4 [3]));
 sky130_fd_sc_hd__nor2_1 \v0/z4/z5/_45_  (.A(\v0/z4/_00_ ),
    .B(\v0/z4/q1 [4]),
    .Y(\v0/z4/z5/_14_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z4/z5/_46_  (.A(\v0/z4/_00_ ),
    .B(\v0/z4/q1 [4]),
    .Y(\v0/z4/z5/_15_ ));
 sky130_fd_sc_hd__nand2b_1 \v0/z4/z5/_47_  (.A_N(\v0/z4/z5/_14_ ),
    .B(\v0/z4/z5/_15_ ),
    .Y(\v0/z4/z5/_16_ ));
 sky130_fd_sc_hd__a21oi_1 \v0/z4/z5/_48_  (.A1(\v0/z4/z5/_10_ ),
    .A2(\v0/z4/z5/_13_ ),
    .B1(\v0/z4/z5/_09_ ),
    .Y(\v0/z4/z5/_17_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z4/z5/_49_  (.A(\v0/z4/z5/_16_ ),
    .B(\v0/z4/z5/_17_ ),
    .Y(\v0/z4/q4 [4]));
 sky130_fd_sc_hd__a311o_1 \v0/z4/z5/_50_  (.A1(\v0/z4/z5/_06_ ),
    .A2(\v0/z4/z5/_10_ ),
    .A3(\v0/z4/z5/_12_ ),
    .B1(\v0/z4/z5/_14_ ),
    .C1(\v0/z4/z5/_09_ ),
    .X(\v0/z4/z5/_18_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z4/z5/_51_  (.A(\v0/z4/z5/_15_ ),
    .B(\v0/z4/z5/_18_ ),
    .Y(\v0/z4/z5/_19_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z4/z5/_52_  (.A(\v0/z4/_01_ ),
    .B(\v0/z4/q1 [5]),
    .Y(\v0/z4/z5/_20_ ));
 sky130_fd_sc_hd__nor2_1 \v0/z4/z5/_53_  (.A(\v0/z4/_01_ ),
    .B(\v0/z4/q1 [5]),
    .Y(\v0/z4/z5/_21_ ));
 sky130_fd_sc_hd__a31oi_1 \v0/z4/z5/_54_  (.A1(\v0/z4/z5/_15_ ),
    .A2(\v0/z4/z5/_18_ ),
    .A3(\v0/z4/z5/_20_ ),
    .B1(\v0/z4/z5/_21_ ),
    .Y(\v0/z4/z5/_22_ ));
 sky130_fd_sc_hd__a21bo_1 \v0/z4/z5/_55_  (.A1(\v0/z4/z5/_20_ ),
    .A2(\v0/z4/z5/_22_ ),
    .B1_N(\v0/z4/z5/_19_ ),
    .X(\v0/z4/z5/_23_ ));
 sky130_fd_sc_hd__o21ai_0 \v0/z4/z5/_56_  (.A1(\v0/z4/z5/_21_ ),
    .A2(\v0/z4/z5/_22_ ),
    .B1(\v0/z4/z5/_23_ ),
    .Y(\v0/z4/q4 [5]));
 sky130_fd_sc_hd__xnor2_1 \v0/z4/z5/_57_  (.A(\v0/z4/_02_ ),
    .B(\v0/z4/q1 [6]),
    .Y(\v0/z4/z5/_24_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z4/z5/_58_  (.A(\v0/z4/z5/_22_ ),
    .B(\v0/z4/z5/_24_ ),
    .Y(\v0/z4/q4 [6]));
 sky130_fd_sc_hd__xnor2_1 \v0/z4/z5/_59_  (.A(\v0/z4/_03_ ),
    .B(\v0/z4/q1 [7]),
    .Y(\v0/z4/z5/_25_ ));
 sky130_fd_sc_hd__maj3_1 \v0/z4/z5/_60_  (.A(\v0/z4/_02_ ),
    .B(\v0/z4/q1 [6]),
    .C(\v0/z4/z5/_22_ ),
    .X(\v0/z4/z5/_26_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z4/z5/_61_  (.A(\v0/z4/z5/_25_ ),
    .B(\v0/z4/z5/_26_ ),
    .Y(\v0/z4/q4 [7]));
 sky130_fd_sc_hd__maj3_1 \v0/z4/z5/_62_  (.A(\v0/z4/_03_ ),
    .B(\v0/z4/q1 [7]),
    .C(\v0/z4/z5/_26_ ),
    .X(\v0/z4/z5/Cout ));
 sky130_fd_sc_hd__xnor2_1 \v0/z4/z6/_050_  (.A(\v0/z4/_09_ ),
    .B(\v0/z4/q2 [0]),
    .Y(\v0/z4/z6/_000_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z4/z6/_051_  (.A(\v0/z4/_13_ ),
    .B(\v0/z4/z6/_000_ ),
    .Y(\v0/z4/q5 [0]));
 sky130_fd_sc_hd__maj3_1 \v0/z4/z6/_052_  (.A(\v0/z4/_09_ ),
    .B(\v0/z4/q2 [0]),
    .C(\v0/z4/_13_ ),
    .X(\v0/z4/z6/_001_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z4/z6/_053_  (.A(\v0/z4/_10_ ),
    .B(\v0/z4/q2 [1]),
    .Y(\v0/z4/z6/_002_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z4/z6/_054_  (.A(\v0/z4/z6/_001_ ),
    .B(\v0/z4/z6/_002_ ),
    .Y(\v0/z4/q5 [1]));
 sky130_fd_sc_hd__maj3_1 \v0/z4/z6/_055_  (.A(\v0/z4/_10_ ),
    .B(\v0/z4/q2 [1]),
    .C(\v0/z4/z6/_001_ ),
    .X(\v0/z4/z6/_003_ ));
 sky130_fd_sc_hd__lpflow_inputiso1p_1 \v0/z4/z6/_056_  (.A(\v0/z4/_11_ ),
    .SLEEP(\v0/z4/q2 [2]),
    .X(\v0/z4/z6/_004_ ));
 sky130_fd_sc_hd__and2_0 \v0/z4/z6/_057_  (.A(\v0/z4/_11_ ),
    .B(\v0/z4/q2 [2]),
    .X(\v0/z4/z6/_005_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z4/z6/_058_  (.A(\v0/z4/_11_ ),
    .B(\v0/z4/q2 [2]),
    .Y(\v0/z4/z6/_006_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z4/z6/_059_  (.A(\v0/z4/z6/_004_ ),
    .B(\v0/z4/z6/_006_ ),
    .Y(\v0/z4/z6/_007_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z4/z6/_060_  (.A(\v0/z4/z6/_003_ ),
    .B(\v0/z4/z6/_007_ ),
    .Y(\v0/z4/q5 [2]));
 sky130_fd_sc_hd__nor2_1 \v0/z4/z6/_061_  (.A(\v0/z4/_12_ ),
    .B(\v0/z4/q2 [3]),
    .Y(\v0/z4/z6/_008_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z4/z6/_062_  (.A(\v0/z4/_12_ ),
    .B(\v0/z4/q2 [3]),
    .Y(\v0/z4/z6/_009_ ));
 sky130_fd_sc_hd__clkinv_1 \v0/z4/z6/_063_  (.A(\v0/z4/z6/_009_ ),
    .Y(\v0/z4/z6/_010_ ));
 sky130_fd_sc_hd__nor2_1 \v0/z4/z6/_064_  (.A(\v0/z4/z6/_008_ ),
    .B(\v0/z4/z6/_010_ ),
    .Y(\v0/z4/z6/_011_ ));
 sky130_fd_sc_hd__o21ai_0 \v0/z4/z6/_065_  (.A1(\v0/z4/z6/_003_ ),
    .A2(\v0/z4/z6/_005_ ),
    .B1(\v0/z4/z6/_004_ ),
    .Y(\v0/z4/z6/_012_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z4/z6/_066_  (.A(\v0/z4/z6/_011_ ),
    .B(\v0/z4/z6/_012_ ),
    .Y(\v0/z4/q5 [3]));
 sky130_fd_sc_hd__lpflow_inputiso1p_1 \v0/z4/z6/_067_  (.A(\v0/z4/q3 [0]),
    .SLEEP(\v0/z4/q2 [4]),
    .X(\v0/z4/z6/_013_ ));
 sky130_fd_sc_hd__and2_0 \v0/z4/z6/_068_  (.A(\v0/z4/q3 [0]),
    .B(\v0/z4/q2 [4]),
    .X(\v0/z4/z6/_014_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z4/z6/_069_  (.A(\v0/z4/q3 [0]),
    .B(\v0/z4/q2 [4]),
    .Y(\v0/z4/z6/_015_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z4/z6/_070_  (.A(\v0/z4/z6/_013_ ),
    .B(\v0/z4/z6/_015_ ),
    .Y(\v0/z4/z6/_016_ ));
 sky130_fd_sc_hd__o221a_1 \v0/z4/z6/_071_  (.A1(\v0/z4/_12_ ),
    .A2(\v0/z4/q2 [3]),
    .B1(\v0/z4/z6/_003_ ),
    .B2(\v0/z4/z6/_005_ ),
    .C1(\v0/z4/z6/_004_ ),
    .X(\v0/z4/z6/_017_ ));
 sky130_fd_sc_hd__a21oi_1 \v0/z4/z6/_072_  (.A1(\v0/z4/z6/_009_ ),
    .A2(\v0/z4/z6/_012_ ),
    .B1(\v0/z4/z6/_008_ ),
    .Y(\v0/z4/z6/_018_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z4/z6/_073_  (.A(\v0/z4/z6/_016_ ),
    .B(\v0/z4/z6/_018_ ),
    .Y(\v0/z4/q5 [4]));
 sky130_fd_sc_hd__lpflow_inputiso1p_1 \v0/z4/z6/_074_  (.A(\v0/z4/q3 [1]),
    .SLEEP(\v0/z4/q2 [5]),
    .X(\v0/z4/z6/_019_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z4/z6/_075_  (.A(\v0/z4/q3 [1]),
    .B(\v0/z4/q2 [5]),
    .Y(\v0/z4/z6/_020_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z4/z6/_076_  (.A(\v0/z4/z6/_019_ ),
    .B(\v0/z4/z6/_020_ ),
    .Y(\v0/z4/z6/_021_ ));
 sky130_fd_sc_hd__o21ai_0 \v0/z4/z6/_077_  (.A1(\v0/z4/z6/_014_ ),
    .A2(\v0/z4/z6/_018_ ),
    .B1(\v0/z4/z6/_013_ ),
    .Y(\v0/z4/z6/_022_ ));
 sky130_fd_sc_hd__xor2_1 \v0/z4/z6/_078_  (.A(\v0/z4/z6/_021_ ),
    .B(\v0/z4/z6/_022_ ),
    .X(\v0/z4/q5 [5]));
 sky130_fd_sc_hd__nor2_1 \v0/z4/z6/_079_  (.A(\v0/z4/q3 [2]),
    .B(\v0/z4/q2 [6]),
    .Y(\v0/z4/z6/_023_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z4/z6/_080_  (.A(\v0/z4/q3 [2]),
    .B(\v0/z4/q2 [6]),
    .Y(\v0/z4/z6/_024_ ));
 sky130_fd_sc_hd__nor2b_1 \v0/z4/z6/_081_  (.A(\v0/z4/z6/_023_ ),
    .B_N(\v0/z4/z6/_024_ ),
    .Y(\v0/z4/z6/_025_ ));
 sky130_fd_sc_hd__o311ai_0 \v0/z4/z6/_082_  (.A1(\v0/z4/z6/_010_ ),
    .A2(\v0/z4/z6/_014_ ),
    .A3(\v0/z4/z6/_017_ ),
    .B1(\v0/z4/z6/_019_ ),
    .C1(\v0/z4/z6/_013_ ),
    .Y(\v0/z4/z6/_026_ ));
 sky130_fd_sc_hd__and2_0 \v0/z4/z6/_083_  (.A(\v0/z4/z6/_020_ ),
    .B(\v0/z4/z6/_026_ ),
    .X(\v0/z4/z6/_027_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z4/z6/_084_  (.A(\v0/z4/z6/_025_ ),
    .B(\v0/z4/z6/_027_ ),
    .Y(\v0/z4/q5 [6]));
 sky130_fd_sc_hd__nor2_1 \v0/z4/z6/_085_  (.A(\v0/z4/q3 [3]),
    .B(\v0/z4/q2 [7]),
    .Y(\v0/z4/z6/_028_ ));
 sky130_fd_sc_hd__and2_0 \v0/z4/z6/_086_  (.A(\v0/z4/q3 [3]),
    .B(\v0/z4/q2 [7]),
    .X(\v0/z4/z6/_029_ ));
 sky130_fd_sc_hd__nor2_1 \v0/z4/z6/_087_  (.A(\v0/z4/z6/_028_ ),
    .B(\v0/z4/z6/_029_ ),
    .Y(\v0/z4/z6/_030_ ));
 sky130_fd_sc_hd__a21oi_1 \v0/z4/z6/_088_  (.A1(\v0/z4/z6/_024_ ),
    .A2(\v0/z4/z6/_027_ ),
    .B1(\v0/z4/z6/_023_ ),
    .Y(\v0/z4/z6/_031_ ));
 sky130_fd_sc_hd__xor2_1 \v0/z4/z6/_089_  (.A(\v0/z4/z6/_030_ ),
    .B(\v0/z4/z6/_031_ ),
    .X(\v0/z4/q5 [7]));
 sky130_fd_sc_hd__lpflow_inputiso1p_1 \v0/z4/z6/_090_  (.A(\v0/z4/q3 [4]),
    .SLEEP(\v0/z4/_05_ ),
    .X(\v0/z4/z6/_032_ ));
 sky130_fd_sc_hd__and2_0 \v0/z4/z6/_091_  (.A(\v0/z4/q3 [4]),
    .B(\v0/z4/_05_ ),
    .X(\v0/z4/z6/_033_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z4/z6/_092_  (.A(\v0/z4/q3 [4]),
    .B(\v0/z4/_05_ ),
    .Y(\v0/z4/z6/_034_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z4/z6/_093_  (.A(\v0/z4/z6/_032_ ),
    .B(\v0/z4/z6/_034_ ),
    .Y(\v0/z4/z6/_035_ ));
 sky130_fd_sc_hd__a311oi_1 \v0/z4/z6/_094_  (.A1(\v0/z4/z6/_020_ ),
    .A2(\v0/z4/z6/_024_ ),
    .A3(\v0/z4/z6/_026_ ),
    .B1(\v0/z4/z6/_028_ ),
    .C1(\v0/z4/z6/_023_ ),
    .Y(\v0/z4/z6/_036_ ));
 sky130_fd_sc_hd__lpflow_inputiso1p_1 \v0/z4/z6/_095_  (.A(\v0/z4/z6/_029_ ),
    .SLEEP(\v0/z4/z6/_036_ ),
    .X(\v0/z4/z6/_037_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z4/z6/_096_  (.A(\v0/z4/z6/_035_ ),
    .B(\v0/z4/z6/_037_ ),
    .Y(\v0/z4/q5 [8]));
 sky130_fd_sc_hd__lpflow_inputiso1p_1 \v0/z4/z6/_097_  (.A(\v0/z4/q3 [5]),
    .SLEEP(\v0/z4/_06_ ),
    .X(\v0/z4/z6/_038_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z4/z6/_098_  (.A(\v0/z4/q3 [5]),
    .B(\v0/z4/_06_ ),
    .Y(\v0/z4/z6/_039_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z4/z6/_099_  (.A(\v0/z4/z6/_038_ ),
    .B(\v0/z4/z6/_039_ ),
    .Y(\v0/z4/z6/_040_ ));
 sky130_fd_sc_hd__o21ai_0 \v0/z4/z6/_100_  (.A1(\v0/z4/z6/_033_ ),
    .A2(\v0/z4/z6/_037_ ),
    .B1(\v0/z4/z6/_032_ ),
    .Y(\v0/z4/z6/_041_ ));
 sky130_fd_sc_hd__xor2_1 \v0/z4/z6/_101_  (.A(\v0/z4/z6/_040_ ),
    .B(\v0/z4/z6/_041_ ),
    .X(\v0/z4/q5 [9]));
 sky130_fd_sc_hd__nor2_1 \v0/z4/z6/_102_  (.A(\v0/z4/q3 [6]),
    .B(\v0/z4/_07_ ),
    .Y(\v0/z4/z6/_042_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z4/z6/_103_  (.A(\v0/z4/q3 [6]),
    .B(\v0/z4/_07_ ),
    .Y(\v0/z4/z6/_043_ ));
 sky130_fd_sc_hd__nand2b_1 \v0/z4/z6/_104_  (.A_N(\v0/z4/z6/_042_ ),
    .B(\v0/z4/z6/_043_ ),
    .Y(\v0/z4/z6/_044_ ));
 sky130_fd_sc_hd__o311ai_0 \v0/z4/z6/_105_  (.A1(\v0/z4/z6/_029_ ),
    .A2(\v0/z4/z6/_033_ ),
    .A3(\v0/z4/z6/_036_ ),
    .B1(\v0/z4/z6/_038_ ),
    .C1(\v0/z4/z6/_032_ ),
    .Y(\v0/z4/z6/_045_ ));
 sky130_fd_sc_hd__a21oi_1 \v0/z4/z6/_106_  (.A1(\v0/z4/z6/_039_ ),
    .A2(\v0/z4/z6/_045_ ),
    .B1(\v0/z4/z6/_044_ ),
    .Y(\v0/z4/z6/_046_ ));
 sky130_fd_sc_hd__and3_1 \v0/z4/z6/_107_  (.A(\v0/z4/z6/_039_ ),
    .B(\v0/z4/z6/_044_ ),
    .C(\v0/z4/z6/_045_ ),
    .X(\v0/z4/z6/_047_ ));
 sky130_fd_sc_hd__nor2_1 \v0/z4/z6/_108_  (.A(\v0/z4/z6/_046_ ),
    .B(\v0/z4/z6/_047_ ),
    .Y(\v0/z4/q5 [10]));
 sky130_fd_sc_hd__xnor2_1 \v0/z4/z6/_109_  (.A(\v0/z4/q3 [7]),
    .B(\v0/z4/_08_ ),
    .Y(\v0/z4/z6/_048_ ));
 sky130_fd_sc_hd__a31oi_1 \v0/z4/z6/_110_  (.A1(\v0/z4/z6/_039_ ),
    .A2(\v0/z4/z6/_043_ ),
    .A3(\v0/z4/z6/_045_ ),
    .B1(\v0/z4/z6/_042_ ),
    .Y(\v0/z4/z6/_049_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z4/z6/_111_  (.A(\v0/z4/z6/_048_ ),
    .B(\v0/z4/z6/_049_ ),
    .Y(\v0/z4/q5 [11]));
 sky130_fd_sc_hd__maj3_1 \v0/z4/z6/_112_  (.A(\v0/z4/q3 [7]),
    .B(\v0/z4/_08_ ),
    .C(\v0/z4/z6/_049_ ),
    .X(\v0/z4/z6/Cout ));
 sky130_fd_sc_hd__xnor2_1 \v0/z4/z7/_050_  (.A(\v0/z4/q5 [0]),
    .B(\v0/z4/q4 [0]),
    .Y(\v0/z4/z7/_000_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z4/z7/_051_  (.A(\v0/z4/_18_ ),
    .B(\v0/z4/z7/_000_ ),
    .Y(\v0/q3 [4]));
 sky130_fd_sc_hd__maj3_1 \v0/z4/z7/_052_  (.A(\v0/z4/q5 [0]),
    .B(\v0/z4/q4 [0]),
    .C(\v0/z4/_18_ ),
    .X(\v0/z4/z7/_001_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z4/z7/_053_  (.A(\v0/z4/q5 [1]),
    .B(\v0/z4/q4 [1]),
    .Y(\v0/z4/z7/_002_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z4/z7/_054_  (.A(\v0/z4/z7/_001_ ),
    .B(\v0/z4/z7/_002_ ),
    .Y(\v0/q3 [5]));
 sky130_fd_sc_hd__maj3_1 \v0/z4/z7/_055_  (.A(\v0/z4/q5 [1]),
    .B(\v0/z4/q4 [1]),
    .C(\v0/z4/z7/_001_ ),
    .X(\v0/z4/z7/_003_ ));
 sky130_fd_sc_hd__lpflow_inputiso1p_1 \v0/z4/z7/_056_  (.A(\v0/z4/q5 [2]),
    .SLEEP(\v0/z4/q4 [2]),
    .X(\v0/z4/z7/_004_ ));
 sky130_fd_sc_hd__and2_0 \v0/z4/z7/_057_  (.A(\v0/z4/q5 [2]),
    .B(\v0/z4/q4 [2]),
    .X(\v0/z4/z7/_005_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z4/z7/_058_  (.A(\v0/z4/q5 [2]),
    .B(\v0/z4/q4 [2]),
    .Y(\v0/z4/z7/_006_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z4/z7/_059_  (.A(\v0/z4/z7/_004_ ),
    .B(\v0/z4/z7/_006_ ),
    .Y(\v0/z4/z7/_007_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z4/z7/_060_  (.A(\v0/z4/z7/_003_ ),
    .B(\v0/z4/z7/_007_ ),
    .Y(\v0/q3 [6]));
 sky130_fd_sc_hd__nor2_1 \v0/z4/z7/_061_  (.A(\v0/z4/q5 [3]),
    .B(\v0/z4/q4 [3]),
    .Y(\v0/z4/z7/_008_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z4/z7/_062_  (.A(\v0/z4/q5 [3]),
    .B(\v0/z4/q4 [3]),
    .Y(\v0/z4/z7/_009_ ));
 sky130_fd_sc_hd__clkinv_1 \v0/z4/z7/_063_  (.A(\v0/z4/z7/_009_ ),
    .Y(\v0/z4/z7/_010_ ));
 sky130_fd_sc_hd__nor2_1 \v0/z4/z7/_064_  (.A(\v0/z4/z7/_008_ ),
    .B(\v0/z4/z7/_010_ ),
    .Y(\v0/z4/z7/_011_ ));
 sky130_fd_sc_hd__o21ai_0 \v0/z4/z7/_065_  (.A1(\v0/z4/z7/_003_ ),
    .A2(\v0/z4/z7/_005_ ),
    .B1(\v0/z4/z7/_004_ ),
    .Y(\v0/z4/z7/_012_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z4/z7/_066_  (.A(\v0/z4/z7/_011_ ),
    .B(\v0/z4/z7/_012_ ),
    .Y(\v0/q3 [7]));
 sky130_fd_sc_hd__lpflow_inputiso1p_1 \v0/z4/z7/_067_  (.A(\v0/z4/q5 [4]),
    .SLEEP(\v0/z4/q4 [4]),
    .X(\v0/z4/z7/_013_ ));
 sky130_fd_sc_hd__and2_0 \v0/z4/z7/_068_  (.A(\v0/z4/q5 [4]),
    .B(\v0/z4/q4 [4]),
    .X(\v0/z4/z7/_014_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z4/z7/_069_  (.A(\v0/z4/q5 [4]),
    .B(\v0/z4/q4 [4]),
    .Y(\v0/z4/z7/_015_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z4/z7/_070_  (.A(\v0/z4/z7/_013_ ),
    .B(\v0/z4/z7/_015_ ),
    .Y(\v0/z4/z7/_016_ ));
 sky130_fd_sc_hd__o221a_1 \v0/z4/z7/_071_  (.A1(\v0/z4/q5 [3]),
    .A2(\v0/z4/q4 [3]),
    .B1(\v0/z4/z7/_003_ ),
    .B2(\v0/z4/z7/_005_ ),
    .C1(\v0/z4/z7/_004_ ),
    .X(\v0/z4/z7/_017_ ));
 sky130_fd_sc_hd__a21oi_1 \v0/z4/z7/_072_  (.A1(\v0/z4/z7/_009_ ),
    .A2(\v0/z4/z7/_012_ ),
    .B1(\v0/z4/z7/_008_ ),
    .Y(\v0/z4/z7/_018_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z4/z7/_073_  (.A(\v0/z4/z7/_016_ ),
    .B(\v0/z4/z7/_018_ ),
    .Y(\v0/q3 [8]));
 sky130_fd_sc_hd__lpflow_inputiso1p_1 \v0/z4/z7/_074_  (.A(\v0/z4/q5 [5]),
    .SLEEP(\v0/z4/q4 [5]),
    .X(\v0/z4/z7/_019_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z4/z7/_075_  (.A(\v0/z4/q5 [5]),
    .B(\v0/z4/q4 [5]),
    .Y(\v0/z4/z7/_020_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z4/z7/_076_  (.A(\v0/z4/z7/_019_ ),
    .B(\v0/z4/z7/_020_ ),
    .Y(\v0/z4/z7/_021_ ));
 sky130_fd_sc_hd__o21ai_0 \v0/z4/z7/_077_  (.A1(\v0/z4/z7/_014_ ),
    .A2(\v0/z4/z7/_018_ ),
    .B1(\v0/z4/z7/_013_ ),
    .Y(\v0/z4/z7/_022_ ));
 sky130_fd_sc_hd__xor2_1 \v0/z4/z7/_078_  (.A(\v0/z4/z7/_021_ ),
    .B(\v0/z4/z7/_022_ ),
    .X(\v0/q3 [9]));
 sky130_fd_sc_hd__nor2_1 \v0/z4/z7/_079_  (.A(\v0/z4/q5 [6]),
    .B(\v0/z4/q4 [6]),
    .Y(\v0/z4/z7/_023_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z4/z7/_080_  (.A(\v0/z4/q5 [6]),
    .B(\v0/z4/q4 [6]),
    .Y(\v0/z4/z7/_024_ ));
 sky130_fd_sc_hd__nor2b_1 \v0/z4/z7/_081_  (.A(\v0/z4/z7/_023_ ),
    .B_N(\v0/z4/z7/_024_ ),
    .Y(\v0/z4/z7/_025_ ));
 sky130_fd_sc_hd__o311ai_0 \v0/z4/z7/_082_  (.A1(\v0/z4/z7/_010_ ),
    .A2(\v0/z4/z7/_014_ ),
    .A3(\v0/z4/z7/_017_ ),
    .B1(\v0/z4/z7/_019_ ),
    .C1(\v0/z4/z7/_013_ ),
    .Y(\v0/z4/z7/_026_ ));
 sky130_fd_sc_hd__and2_0 \v0/z4/z7/_083_  (.A(\v0/z4/z7/_020_ ),
    .B(\v0/z4/z7/_026_ ),
    .X(\v0/z4/z7/_027_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z4/z7/_084_  (.A(\v0/z4/z7/_025_ ),
    .B(\v0/z4/z7/_027_ ),
    .Y(\v0/q3 [10]));
 sky130_fd_sc_hd__nor2_1 \v0/z4/z7/_085_  (.A(\v0/z4/q5 [7]),
    .B(\v0/z4/q4 [7]),
    .Y(\v0/z4/z7/_028_ ));
 sky130_fd_sc_hd__and2_0 \v0/z4/z7/_086_  (.A(\v0/z4/q5 [7]),
    .B(\v0/z4/q4 [7]),
    .X(\v0/z4/z7/_029_ ));
 sky130_fd_sc_hd__nor2_1 \v0/z4/z7/_087_  (.A(\v0/z4/z7/_028_ ),
    .B(\v0/z4/z7/_029_ ),
    .Y(\v0/z4/z7/_030_ ));
 sky130_fd_sc_hd__a21oi_1 \v0/z4/z7/_088_  (.A1(\v0/z4/z7/_024_ ),
    .A2(\v0/z4/z7/_027_ ),
    .B1(\v0/z4/z7/_023_ ),
    .Y(\v0/z4/z7/_031_ ));
 sky130_fd_sc_hd__xor2_1 \v0/z4/z7/_089_  (.A(\v0/z4/z7/_030_ ),
    .B(\v0/z4/z7/_031_ ),
    .X(\v0/q3 [11]));
 sky130_fd_sc_hd__lpflow_inputiso1p_1 \v0/z4/z7/_090_  (.A(\v0/z4/q5 [8]),
    .SLEEP(\v0/z4/_14_ ),
    .X(\v0/z4/z7/_032_ ));
 sky130_fd_sc_hd__and2_0 \v0/z4/z7/_091_  (.A(\v0/z4/q5 [8]),
    .B(\v0/z4/_14_ ),
    .X(\v0/z4/z7/_033_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z4/z7/_092_  (.A(\v0/z4/q5 [8]),
    .B(\v0/z4/_14_ ),
    .Y(\v0/z4/z7/_034_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z4/z7/_093_  (.A(\v0/z4/z7/_032_ ),
    .B(\v0/z4/z7/_034_ ),
    .Y(\v0/z4/z7/_035_ ));
 sky130_fd_sc_hd__a311oi_1 \v0/z4/z7/_094_  (.A1(\v0/z4/z7/_020_ ),
    .A2(\v0/z4/z7/_024_ ),
    .A3(\v0/z4/z7/_026_ ),
    .B1(\v0/z4/z7/_028_ ),
    .C1(\v0/z4/z7/_023_ ),
    .Y(\v0/z4/z7/_036_ ));
 sky130_fd_sc_hd__lpflow_inputiso1p_1 \v0/z4/z7/_095_  (.A(\v0/z4/z7/_029_ ),
    .SLEEP(\v0/z4/z7/_036_ ),
    .X(\v0/z4/z7/_037_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z4/z7/_096_  (.A(\v0/z4/z7/_035_ ),
    .B(\v0/z4/z7/_037_ ),
    .Y(\v0/q3 [12]));
 sky130_fd_sc_hd__lpflow_inputiso1p_1 \v0/z4/z7/_097_  (.A(\v0/z4/q5 [9]),
    .SLEEP(\v0/z4/_15_ ),
    .X(\v0/z4/z7/_038_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z4/z7/_098_  (.A(\v0/z4/q5 [9]),
    .B(\v0/z4/_15_ ),
    .Y(\v0/z4/z7/_039_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z4/z7/_099_  (.A(\v0/z4/z7/_038_ ),
    .B(\v0/z4/z7/_039_ ),
    .Y(\v0/z4/z7/_040_ ));
 sky130_fd_sc_hd__o21ai_0 \v0/z4/z7/_100_  (.A1(\v0/z4/z7/_033_ ),
    .A2(\v0/z4/z7/_037_ ),
    .B1(\v0/z4/z7/_032_ ),
    .Y(\v0/z4/z7/_041_ ));
 sky130_fd_sc_hd__xor2_1 \v0/z4/z7/_101_  (.A(\v0/z4/z7/_040_ ),
    .B(\v0/z4/z7/_041_ ),
    .X(\v0/q3 [13]));
 sky130_fd_sc_hd__nor2_1 \v0/z4/z7/_102_  (.A(\v0/z4/q5 [10]),
    .B(\v0/z4/_16_ ),
    .Y(\v0/z4/z7/_042_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z4/z7/_103_  (.A(\v0/z4/q5 [10]),
    .B(\v0/z4/_16_ ),
    .Y(\v0/z4/z7/_043_ ));
 sky130_fd_sc_hd__nand2b_1 \v0/z4/z7/_104_  (.A_N(\v0/z4/z7/_042_ ),
    .B(\v0/z4/z7/_043_ ),
    .Y(\v0/z4/z7/_044_ ));
 sky130_fd_sc_hd__o311ai_0 \v0/z4/z7/_105_  (.A1(\v0/z4/z7/_029_ ),
    .A2(\v0/z4/z7/_033_ ),
    .A3(\v0/z4/z7/_036_ ),
    .B1(\v0/z4/z7/_038_ ),
    .C1(\v0/z4/z7/_032_ ),
    .Y(\v0/z4/z7/_045_ ));
 sky130_fd_sc_hd__a21oi_1 \v0/z4/z7/_106_  (.A1(\v0/z4/z7/_039_ ),
    .A2(\v0/z4/z7/_045_ ),
    .B1(\v0/z4/z7/_044_ ),
    .Y(\v0/z4/z7/_046_ ));
 sky130_fd_sc_hd__and3_1 \v0/z4/z7/_107_  (.A(\v0/z4/z7/_039_ ),
    .B(\v0/z4/z7/_044_ ),
    .C(\v0/z4/z7/_045_ ),
    .X(\v0/z4/z7/_047_ ));
 sky130_fd_sc_hd__nor2_1 \v0/z4/z7/_108_  (.A(\v0/z4/z7/_046_ ),
    .B(\v0/z4/z7/_047_ ),
    .Y(\v0/q3 [14]));
 sky130_fd_sc_hd__xnor2_1 \v0/z4/z7/_109_  (.A(\v0/z4/q5 [11]),
    .B(\v0/z4/_17_ ),
    .Y(\v0/z4/z7/_048_ ));
 sky130_fd_sc_hd__a31oi_1 \v0/z4/z7/_110_  (.A1(\v0/z4/z7/_039_ ),
    .A2(\v0/z4/z7/_043_ ),
    .A3(\v0/z4/z7/_045_ ),
    .B1(\v0/z4/z7/_042_ ),
    .Y(\v0/z4/z7/_049_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z4/z7/_111_  (.A(\v0/z4/z7/_048_ ),
    .B(\v0/z4/z7/_049_ ),
    .Y(\v0/q3 [15]));
 sky130_fd_sc_hd__maj3_1 \v0/z4/z7/_112_  (.A(\v0/z4/q5 [11]),
    .B(\v0/z4/_17_ ),
    .C(\v0/z4/z7/_049_ ),
    .X(\v0/z4/z7/Cout ));
 sky130_fd_sc_hd__xnor2_1 \v0/z5/_070_  (.A(\v0/q0 [8]),
    .B(\v0/q1 [0]),
    .Y(\v0/z5/_030_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z5/_071_  (.A(\v0/_08_ ),
    .B(\v0/z5/_030_ ),
    .Y(\v0/q4 [0]));
 sky130_fd_sc_hd__maj3_1 \v0/z5/_072_  (.A(\v0/q0 [8]),
    .B(\v0/q1 [0]),
    .C(\v0/_08_ ),
    .X(\v0/z5/_031_ ));
 sky130_fd_sc_hd__lpflow_inputiso1p_1 \v0/z5/_073_  (.A(\v0/q0 [9]),
    .SLEEP(\v0/q1 [1]),
    .X(\v0/z5/_032_ ));
 sky130_fd_sc_hd__and2_0 \v0/z5/_074_  (.A(\v0/q0 [9]),
    .B(\v0/q1 [1]),
    .X(\v0/z5/_033_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z5/_075_  (.A(\v0/q0 [9]),
    .B(\v0/q1 [1]),
    .Y(\v0/z5/_034_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z5/_076_  (.A(\v0/z5/_032_ ),
    .B(\v0/z5/_034_ ),
    .Y(\v0/z5/_035_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z5/_077_  (.A(\v0/z5/_031_ ),
    .B(\v0/z5/_035_ ),
    .Y(\v0/q4 [1]));
 sky130_fd_sc_hd__nand2_1 \v0/z5/_078_  (.A(\v0/q0 [10]),
    .B(\v0/q1 [2]),
    .Y(\v0/z5/_036_ ));
 sky130_fd_sc_hd__xor2_1 \v0/z5/_079_  (.A(\v0/q0 [10]),
    .B(\v0/q1 [2]),
    .X(\v0/z5/_037_ ));
 sky130_fd_sc_hd__o21ai_0 \v0/z5/_080_  (.A1(\v0/z5/_031_ ),
    .A2(\v0/z5/_033_ ),
    .B1(\v0/z5/_032_ ),
    .Y(\v0/z5/_038_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z5/_081_  (.A(\v0/z5/_037_ ),
    .B(\v0/z5/_038_ ),
    .Y(\v0/q4 [2]));
 sky130_fd_sc_hd__nor2_1 \v0/z5/_082_  (.A(\v0/q0 [11]),
    .B(\v0/q1 [3]),
    .Y(\v0/z5/_039_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z5/_083_  (.A(\v0/q0 [11]),
    .B(\v0/q1 [3]),
    .Y(\v0/z5/_040_ ));
 sky130_fd_sc_hd__nand2b_1 \v0/z5/_084_  (.A_N(\v0/z5/_039_ ),
    .B(\v0/z5/_040_ ),
    .Y(\v0/z5/_041_ ));
 sky130_fd_sc_hd__o221ai_1 \v0/z5/_085_  (.A1(\v0/q0 [10]),
    .A2(\v0/q1 [2]),
    .B1(\v0/z5/_031_ ),
    .B2(\v0/z5/_033_ ),
    .C1(\v0/z5/_032_ ),
    .Y(\v0/z5/_042_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z5/_086_  (.A(\v0/z5/_036_ ),
    .B(\v0/z5/_042_ ),
    .Y(\v0/z5/_043_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z5/_087_  (.A(\v0/z5/_041_ ),
    .B(\v0/z5/_043_ ),
    .Y(\v0/q4 [3]));
 sky130_fd_sc_hd__nand2_1 \v0/z5/_088_  (.A(\v0/q0 [12]),
    .B(\v0/q1 [4]),
    .Y(\v0/z5/_044_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z5/_089_  (.A(\v0/q0 [12]),
    .B(\v0/q1 [4]),
    .Y(\v0/z5/_045_ ));
 sky130_fd_sc_hd__a31oi_1 \v0/z5/_090_  (.A1(\v0/z5/_036_ ),
    .A2(\v0/z5/_040_ ),
    .A3(\v0/z5/_042_ ),
    .B1(\v0/z5/_039_ ),
    .Y(\v0/z5/_046_ ));
 sky130_fd_sc_hd__a311oi_1 \v0/z5/_091_  (.A1(\v0/z5/_036_ ),
    .A2(\v0/z5/_040_ ),
    .A3(\v0/z5/_042_ ),
    .B1(\v0/z5/_045_ ),
    .C1(\v0/z5/_039_ ),
    .Y(\v0/z5/_047_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z5/_092_  (.A(\v0/z5/_045_ ),
    .B(\v0/z5/_046_ ),
    .Y(\v0/q4 [4]));
 sky130_fd_sc_hd__nor2_1 \v0/z5/_093_  (.A(\v0/q0 [13]),
    .B(\v0/q1 [5]),
    .Y(\v0/z5/_048_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z5/_094_  (.A(\v0/q0 [13]),
    .B(\v0/q1 [5]),
    .Y(\v0/z5/_049_ ));
 sky130_fd_sc_hd__nor2b_1 \v0/z5/_095_  (.A(\v0/z5/_048_ ),
    .B_N(\v0/z5/_049_ ),
    .Y(\v0/z5/_050_ ));
 sky130_fd_sc_hd__a21oi_1 \v0/z5/_096_  (.A1(\v0/q0 [12]),
    .A2(\v0/q1 [4]),
    .B1(\v0/z5/_047_ ),
    .Y(\v0/z5/_051_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z5/_097_  (.A(\v0/z5/_050_ ),
    .B(\v0/z5/_051_ ),
    .Y(\v0/q4 [5]));
 sky130_fd_sc_hd__nand2_1 \v0/z5/_098_  (.A(\v0/q0 [14]),
    .B(\v0/q1 [6]),
    .Y(\v0/z5/_052_ ));
 sky130_fd_sc_hd__xor2_1 \v0/z5/_099_  (.A(\v0/q0 [14]),
    .B(\v0/q1 [6]),
    .X(\v0/z5/_053_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z5/_100_  (.A(\v0/z5/_044_ ),
    .B(\v0/z5/_049_ ),
    .Y(\v0/z5/_054_ ));
 sky130_fd_sc_hd__o21ai_0 \v0/z5/_101_  (.A1(\v0/z5/_048_ ),
    .A2(\v0/z5/_051_ ),
    .B1(\v0/z5/_049_ ),
    .Y(\v0/z5/_055_ ));
 sky130_fd_sc_hd__o221ai_1 \v0/z5/_102_  (.A1(\v0/q0 [13]),
    .A2(\v0/q1 [5]),
    .B1(\v0/z5/_047_ ),
    .B2(\v0/z5/_054_ ),
    .C1(\v0/z5/_053_ ),
    .Y(\v0/z5/_056_ ));
 sky130_fd_sc_hd__xor2_1 \v0/z5/_103_  (.A(\v0/z5/_053_ ),
    .B(\v0/z5/_055_ ),
    .X(\v0/q4 [6]));
 sky130_fd_sc_hd__nor2_1 \v0/z5/_104_  (.A(\v0/q0 [15]),
    .B(\v0/q1 [7]),
    .Y(\v0/z5/_057_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z5/_105_  (.A(\v0/q0 [15]),
    .B(\v0/q1 [7]),
    .Y(\v0/z5/_058_ ));
 sky130_fd_sc_hd__nor2b_1 \v0/z5/_106_  (.A(\v0/z5/_057_ ),
    .B_N(\v0/z5/_058_ ),
    .Y(\v0/z5/_059_ ));
 sky130_fd_sc_hd__o211ai_1 \v0/z5/_107_  (.A1(\v0/z5/_048_ ),
    .A2(\v0/z5/_051_ ),
    .B1(\v0/z5/_052_ ),
    .C1(\v0/z5/_049_ ),
    .Y(\v0/z5/_060_ ));
 sky130_fd_sc_hd__o21ai_0 \v0/z5/_108_  (.A1(\v0/q0 [14]),
    .A2(\v0/q1 [6]),
    .B1(\v0/z5/_060_ ),
    .Y(\v0/z5/_061_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z5/_109_  (.A(\v0/z5/_059_ ),
    .B(\v0/z5/_061_ ),
    .Y(\v0/q4 [7]));
 sky130_fd_sc_hd__and2_0 \v0/z5/_110_  (.A(\v0/_00_ ),
    .B(\v0/q1 [8]),
    .X(\v0/z5/_062_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z5/_111_  (.A(\v0/_00_ ),
    .B(\v0/q1 [8]),
    .Y(\v0/z5/_063_ ));
 sky130_fd_sc_hd__a31oi_1 \v0/z5/_112_  (.A1(\v0/z5/_052_ ),
    .A2(\v0/z5/_056_ ),
    .A3(\v0/z5/_058_ ),
    .B1(\v0/z5/_057_ ),
    .Y(\v0/z5/_064_ ));
 sky130_fd_sc_hd__a311oi_1 \v0/z5/_113_  (.A1(\v0/z5/_052_ ),
    .A2(\v0/z5/_056_ ),
    .A3(\v0/z5/_058_ ),
    .B1(\v0/z5/_063_ ),
    .C1(\v0/z5/_057_ ),
    .Y(\v0/z5/_065_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z5/_114_  (.A(\v0/z5/_063_ ),
    .B(\v0/z5/_064_ ),
    .Y(\v0/q4 [8]));
 sky130_fd_sc_hd__nand2_1 \v0/z5/_115_  (.A(\v0/_01_ ),
    .B(\v0/q1 [9]),
    .Y(\v0/z5/_066_ ));
 sky130_fd_sc_hd__xor2_1 \v0/z5/_116_  (.A(\v0/_01_ ),
    .B(\v0/q1 [9]),
    .X(\v0/z5/_067_ ));
 sky130_fd_sc_hd__o21ai_0 \v0/z5/_117_  (.A1(\v0/z5/_062_ ),
    .A2(\v0/z5/_065_ ),
    .B1(\v0/z5/_067_ ),
    .Y(\v0/z5/_068_ ));
 sky130_fd_sc_hd__nor3_1 \v0/z5/_118_  (.A(\v0/z5/_062_ ),
    .B(\v0/z5/_065_ ),
    .C(\v0/z5/_067_ ),
    .Y(\v0/z5/_069_ ));
 sky130_fd_sc_hd__lpflow_isobufsrc_1 \v0/z5/_119_  (.A(\v0/z5/_068_ ),
    .SLEEP(\v0/z5/_069_ ),
    .X(\v0/q4 [9]));
 sky130_fd_sc_hd__nor2_1 \v0/z5/_120_  (.A(\v0/_02_ ),
    .B(\v0/q1 [10]),
    .Y(\v0/z5/_000_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z5/_121_  (.A(\v0/_02_ ),
    .B(\v0/q1 [10]),
    .Y(\v0/z5/_001_ ));
 sky130_fd_sc_hd__nand2b_1 \v0/z5/_122_  (.A_N(\v0/z5/_000_ ),
    .B(\v0/z5/_001_ ),
    .Y(\v0/z5/_002_ ));
 sky130_fd_sc_hd__o22ai_1 \v0/z5/_123_  (.A1(\v0/_01_ ),
    .A2(\v0/q1 [9]),
    .B1(\v0/z5/_062_ ),
    .B2(\v0/z5/_065_ ),
    .Y(\v0/z5/_003_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z5/_124_  (.A(\v0/z5/_066_ ),
    .B(\v0/z5/_003_ ),
    .Y(\v0/z5/_004_ ));
 sky130_fd_sc_hd__a21o_1 \v0/z5/_125_  (.A1(\v0/z5/_066_ ),
    .A2(\v0/z5/_003_ ),
    .B1(\v0/z5/_002_ ),
    .X(\v0/z5/_005_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z5/_126_  (.A(\v0/z5/_002_ ),
    .B(\v0/z5/_004_ ),
    .Y(\v0/q4 [10]));
 sky130_fd_sc_hd__nor2_1 \v0/z5/_127_  (.A(\v0/_03_ ),
    .B(\v0/q1 [11]),
    .Y(\v0/z5/_006_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z5/_128_  (.A(\v0/_03_ ),
    .B(\v0/q1 [11]),
    .Y(\v0/z5/_007_ ));
 sky130_fd_sc_hd__nand2b_1 \v0/z5/_129_  (.A_N(\v0/z5/_006_ ),
    .B(\v0/z5/_007_ ),
    .Y(\v0/z5/_008_ ));
 sky130_fd_sc_hd__a31oi_1 \v0/z5/_130_  (.A1(\v0/z5/_066_ ),
    .A2(\v0/z5/_068_ ),
    .A3(\v0/z5/_001_ ),
    .B1(\v0/z5/_000_ ),
    .Y(\v0/z5/_009_ ));
 sky130_fd_sc_hd__a311o_1 \v0/z5/_131_  (.A1(\v0/z5/_066_ ),
    .A2(\v0/z5/_068_ ),
    .A3(\v0/z5/_001_ ),
    .B1(\v0/z5/_008_ ),
    .C1(\v0/z5/_000_ ),
    .X(\v0/z5/_010_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z5/_132_  (.A(\v0/z5/_008_ ),
    .B(\v0/z5/_009_ ),
    .Y(\v0/q4 [11]));
 sky130_fd_sc_hd__nor2_1 \v0/z5/_133_  (.A(\v0/_04_ ),
    .B(\v0/q1 [12]),
    .Y(\v0/z5/_011_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z5/_134_  (.A(\v0/_04_ ),
    .B(\v0/q1 [12]),
    .Y(\v0/z5/_012_ ));
 sky130_fd_sc_hd__nand2b_1 \v0/z5/_135_  (.A_N(\v0/z5/_011_ ),
    .B(\v0/z5/_012_ ),
    .Y(\v0/z5/_013_ ));
 sky130_fd_sc_hd__a31oi_1 \v0/z5/_136_  (.A1(\v0/z5/_001_ ),
    .A2(\v0/z5/_005_ ),
    .A3(\v0/z5/_007_ ),
    .B1(\v0/z5/_006_ ),
    .Y(\v0/z5/_014_ ));
 sky130_fd_sc_hd__a311o_1 \v0/z5/_137_  (.A1(\v0/z5/_001_ ),
    .A2(\v0/z5/_005_ ),
    .A3(\v0/z5/_007_ ),
    .B1(\v0/z5/_013_ ),
    .C1(\v0/z5/_006_ ),
    .X(\v0/z5/_015_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z5/_138_  (.A(\v0/z5/_013_ ),
    .B(\v0/z5/_014_ ),
    .Y(\v0/q4 [12]));
 sky130_fd_sc_hd__nor2_1 \v0/z5/_139_  (.A(\v0/_05_ ),
    .B(\v0/q1 [13]),
    .Y(\v0/z5/_016_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z5/_140_  (.A(\v0/_05_ ),
    .B(\v0/q1 [13]),
    .Y(\v0/z5/_017_ ));
 sky130_fd_sc_hd__nand2b_1 \v0/z5/_141_  (.A_N(\v0/z5/_016_ ),
    .B(\v0/z5/_017_ ),
    .Y(\v0/z5/_018_ ));
 sky130_fd_sc_hd__a31oi_1 \v0/z5/_142_  (.A1(\v0/z5/_007_ ),
    .A2(\v0/z5/_010_ ),
    .A3(\v0/z5/_012_ ),
    .B1(\v0/z5/_011_ ),
    .Y(\v0/z5/_019_ ));
 sky130_fd_sc_hd__a311oi_1 \v0/z5/_143_  (.A1(\v0/z5/_007_ ),
    .A2(\v0/z5/_010_ ),
    .A3(\v0/z5/_012_ ),
    .B1(\v0/z5/_018_ ),
    .C1(\v0/z5/_011_ ),
    .Y(\v0/z5/_020_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z5/_144_  (.A(\v0/z5/_018_ ),
    .B(\v0/z5/_019_ ),
    .Y(\v0/q4 [13]));
 sky130_fd_sc_hd__nand2_1 \v0/z5/_145_  (.A(\v0/_06_ ),
    .B(\v0/q1 [14]),
    .Y(\v0/z5/_021_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z5/_146_  (.A(\v0/_06_ ),
    .B(\v0/q1 [14]),
    .Y(\v0/z5/_022_ ));
 sky130_fd_sc_hd__a31oi_1 \v0/z5/_147_  (.A1(\v0/z5/_012_ ),
    .A2(\v0/z5/_015_ ),
    .A3(\v0/z5/_017_ ),
    .B1(\v0/z5/_016_ ),
    .Y(\v0/z5/_023_ ));
 sky130_fd_sc_hd__a311o_1 \v0/z5/_148_  (.A1(\v0/z5/_012_ ),
    .A2(\v0/z5/_015_ ),
    .A3(\v0/z5/_017_ ),
    .B1(\v0/z5/_022_ ),
    .C1(\v0/z5/_016_ ),
    .X(\v0/z5/_024_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z5/_149_  (.A(\v0/z5/_022_ ),
    .B(\v0/z5/_023_ ),
    .Y(\v0/q4 [14]));
 sky130_fd_sc_hd__nor2_1 \v0/z5/_150_  (.A(\v0/_07_ ),
    .B(\v0/q1 [15]),
    .Y(\v0/z5/_025_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z5/_151_  (.A(\v0/_07_ ),
    .B(\v0/q1 [15]),
    .Y(\v0/z5/_026_ ));
 sky130_fd_sc_hd__nor2b_1 \v0/z5/_152_  (.A(\v0/z5/_025_ ),
    .B_N(\v0/z5/_026_ ),
    .Y(\v0/z5/_027_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z5/_153_  (.A(\v0/z5/_017_ ),
    .B(\v0/z5/_021_ ),
    .Y(\v0/z5/_028_ ));
 sky130_fd_sc_hd__o22ai_1 \v0/z5/_154_  (.A1(\v0/_06_ ),
    .A2(\v0/q1 [14]),
    .B1(\v0/z5/_020_ ),
    .B2(\v0/z5/_028_ ),
    .Y(\v0/z5/_029_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z5/_155_  (.A(\v0/z5/_027_ ),
    .B(\v0/z5/_029_ ),
    .Y(\v0/q4 [15]));
 sky130_fd_sc_hd__a31oi_1 \v0/z5/_156_  (.A1(\v0/z5/_021_ ),
    .A2(\v0/z5/_024_ ),
    .A3(\v0/z5/_026_ ),
    .B1(\v0/z5/_025_ ),
    .Y(\v0/z5/Cout ));
 sky130_fd_sc_hd__xnor2_1 \v0/z6/_113_  (.A(\v0/_17_ ),
    .B(\v0/q2 [0]),
    .Y(\v0/z6/_093_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z6/_114_  (.A(\v0/_25_ ),
    .B(\v0/z6/_093_ ),
    .Y(\v0/q5 [0]));
 sky130_fd_sc_hd__maj3_1 \v0/z6/_115_  (.A(\v0/_17_ ),
    .B(\v0/q2 [0]),
    .C(\v0/_25_ ),
    .X(\v0/z6/_094_ ));
 sky130_fd_sc_hd__lpflow_inputiso1p_1 \v0/z6/_116_  (.A(\v0/_18_ ),
    .SLEEP(\v0/q2 [1]),
    .X(\v0/z6/_095_ ));
 sky130_fd_sc_hd__and2_0 \v0/z6/_117_  (.A(\v0/_18_ ),
    .B(\v0/q2 [1]),
    .X(\v0/z6/_096_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z6/_118_  (.A(\v0/_18_ ),
    .B(\v0/q2 [1]),
    .Y(\v0/z6/_097_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z6/_119_  (.A(\v0/z6/_095_ ),
    .B(\v0/z6/_097_ ),
    .Y(\v0/z6/_098_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z6/_120_  (.A(\v0/z6/_094_ ),
    .B(\v0/z6/_098_ ),
    .Y(\v0/q5 [1]));
 sky130_fd_sc_hd__nor2_1 \v0/z6/_121_  (.A(\v0/_19_ ),
    .B(\v0/q2 [2]),
    .Y(\v0/z6/_099_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z6/_122_  (.A(\v0/_19_ ),
    .B(\v0/q2 [2]),
    .Y(\v0/z6/_100_ ));
 sky130_fd_sc_hd__xor2_1 \v0/z6/_123_  (.A(\v0/_19_ ),
    .B(\v0/q2 [2]),
    .X(\v0/z6/_101_ ));
 sky130_fd_sc_hd__o21ai_0 \v0/z6/_124_  (.A1(\v0/z6/_094_ ),
    .A2(\v0/z6/_096_ ),
    .B1(\v0/z6/_095_ ),
    .Y(\v0/z6/_102_ ));
 sky130_fd_sc_hd__o211a_1 \v0/z6/_125_  (.A1(\v0/z6/_094_ ),
    .A2(\v0/z6/_096_ ),
    .B1(\v0/z6/_101_ ),
    .C1(\v0/z6/_095_ ),
    .X(\v0/z6/_103_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z6/_126_  (.A(\v0/z6/_101_ ),
    .B(\v0/z6/_102_ ),
    .Y(\v0/q5 [2]));
 sky130_fd_sc_hd__nand2_1 \v0/z6/_127_  (.A(\v0/_20_ ),
    .B(\v0/q2 [3]),
    .Y(\v0/z6/_104_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z6/_128_  (.A(\v0/_20_ ),
    .B(\v0/q2 [3]),
    .Y(\v0/z6/_105_ ));
 sky130_fd_sc_hd__o21ai_0 \v0/z6/_129_  (.A1(\v0/z6/_099_ ),
    .A2(\v0/z6/_102_ ),
    .B1(\v0/z6/_100_ ),
    .Y(\v0/z6/_106_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z6/_130_  (.A(\v0/z6/_105_ ),
    .B(\v0/z6/_106_ ),
    .Y(\v0/q5 [3]));
 sky130_fd_sc_hd__lpflow_inputiso1p_1 \v0/z6/_131_  (.A(\v0/_21_ ),
    .SLEEP(\v0/q2 [4]),
    .X(\v0/z6/_107_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z6/_132_  (.A(\v0/_21_ ),
    .B(\v0/q2 [4]),
    .Y(\v0/z6/_108_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z6/_133_  (.A(\v0/z6/_107_ ),
    .B(\v0/z6/_108_ ),
    .Y(\v0/z6/_109_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z6/_134_  (.A(\v0/z6/_100_ ),
    .B(\v0/z6/_104_ ),
    .Y(\v0/z6/_110_ ));
 sky130_fd_sc_hd__o22a_1 \v0/z6/_135_  (.A1(\v0/_20_ ),
    .A2(\v0/q2 [3]),
    .B1(\v0/z6/_103_ ),
    .B2(\v0/z6/_110_ ),
    .X(\v0/z6/_111_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z6/_136_  (.A(\v0/z6/_109_ ),
    .B(\v0/z6/_111_ ),
    .Y(\v0/q5 [4]));
 sky130_fd_sc_hd__nor2_1 \v0/z6/_137_  (.A(\v0/_22_ ),
    .B(\v0/q2 [5]),
    .Y(\v0/z6/_112_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z6/_138_  (.A(\v0/_22_ ),
    .B(\v0/q2 [5]),
    .Y(\v0/z6/_000_ ));
 sky130_fd_sc_hd__nand2b_1 \v0/z6/_139_  (.A_N(\v0/z6/_112_ ),
    .B(\v0/z6/_000_ ),
    .Y(\v0/z6/_001_ ));
 sky130_fd_sc_hd__o221ai_1 \v0/z6/_140_  (.A1(\v0/_20_ ),
    .A2(\v0/q2 [3]),
    .B1(\v0/z6/_103_ ),
    .B2(\v0/z6/_110_ ),
    .C1(\v0/z6/_107_ ),
    .Y(\v0/z6/_002_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z6/_141_  (.A(\v0/z6/_108_ ),
    .B(\v0/z6/_002_ ),
    .Y(\v0/z6/_003_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z6/_142_  (.A(\v0/z6/_001_ ),
    .B(\v0/z6/_003_ ),
    .Y(\v0/q5 [5]));
 sky130_fd_sc_hd__nor2_1 \v0/z6/_143_  (.A(\v0/_23_ ),
    .B(\v0/q2 [6]),
    .Y(\v0/z6/_004_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z6/_144_  (.A(\v0/_23_ ),
    .B(\v0/q2 [6]),
    .Y(\v0/z6/_005_ ));
 sky130_fd_sc_hd__nor2b_1 \v0/z6/_145_  (.A(\v0/z6/_004_ ),
    .B_N(\v0/z6/_005_ ),
    .Y(\v0/z6/_006_ ));
 sky130_fd_sc_hd__clkinv_1 \v0/z6/_146_  (.A(\v0/z6/_006_ ),
    .Y(\v0/z6/_007_ ));
 sky130_fd_sc_hd__o21ai_0 \v0/z6/_147_  (.A1(\v0/_22_ ),
    .A2(\v0/q2 [5]),
    .B1(\v0/z6/_003_ ),
    .Y(\v0/z6/_008_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z6/_148_  (.A(\v0/z6/_000_ ),
    .B(\v0/z6/_008_ ),
    .Y(\v0/z6/_009_ ));
 sky130_fd_sc_hd__a311o_1 \v0/z6/_149_  (.A1(\v0/z6/_108_ ),
    .A2(\v0/z6/_000_ ),
    .A3(\v0/z6/_002_ ),
    .B1(\v0/z6/_007_ ),
    .C1(\v0/z6/_112_ ),
    .X(\v0/z6/_010_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z6/_150_  (.A(\v0/z6/_007_ ),
    .B(\v0/z6/_009_ ),
    .Y(\v0/q5 [6]));
 sky130_fd_sc_hd__nor2_1 \v0/z6/_151_  (.A(\v0/_24_ ),
    .B(\v0/q2 [7]),
    .Y(\v0/z6/_011_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z6/_152_  (.A(\v0/_24_ ),
    .B(\v0/q2 [7]),
    .Y(\v0/z6/_012_ ));
 sky130_fd_sc_hd__a31oi_1 \v0/z6/_153_  (.A1(\v0/z6/_000_ ),
    .A2(\v0/z6/_005_ ),
    .A3(\v0/z6/_008_ ),
    .B1(\v0/z6/_004_ ),
    .Y(\v0/z6/_013_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z6/_154_  (.A(\v0/z6/_012_ ),
    .B(\v0/z6/_013_ ),
    .Y(\v0/q5 [7]));
 sky130_fd_sc_hd__nand2_1 \v0/z6/_155_  (.A(\v0/q3 [0]),
    .B(\v0/q2 [8]),
    .Y(\v0/z6/_014_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z6/_156_  (.A(\v0/q3 [0]),
    .B(\v0/q2 [8]),
    .Y(\v0/z6/_015_ ));
 sky130_fd_sc_hd__a22oi_1 \v0/z6/_157_  (.A1(\v0/_23_ ),
    .A2(\v0/q2 [6]),
    .B1(\v0/_24_ ),
    .B2(\v0/q2 [7]),
    .Y(\v0/z6/_016_ ));
 sky130_fd_sc_hd__a21oi_1 \v0/z6/_158_  (.A1(\v0/z6/_010_ ),
    .A2(\v0/z6/_016_ ),
    .B1(\v0/z6/_011_ ),
    .Y(\v0/z6/_017_ ));
 sky130_fd_sc_hd__a211oi_1 \v0/z6/_159_  (.A1(\v0/z6/_010_ ),
    .A2(\v0/z6/_016_ ),
    .B1(\v0/z6/_015_ ),
    .C1(\v0/z6/_011_ ),
    .Y(\v0/z6/_018_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z6/_160_  (.A(\v0/z6/_015_ ),
    .B(\v0/z6/_017_ ),
    .Y(\v0/q5 [8]));
 sky130_fd_sc_hd__lpflow_inputiso1p_1 \v0/z6/_161_  (.A(\v0/q3 [1]),
    .SLEEP(\v0/q2 [9]),
    .X(\v0/z6/_019_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z6/_162_  (.A(\v0/q3 [1]),
    .B(\v0/q2 [9]),
    .Y(\v0/z6/_020_ ));
 sky130_fd_sc_hd__and2_0 \v0/z6/_163_  (.A(\v0/z6/_019_ ),
    .B(\v0/z6/_020_ ),
    .X(\v0/z6/_021_ ));
 sky130_fd_sc_hd__a21oi_1 \v0/z6/_164_  (.A1(\v0/q3 [0]),
    .A2(\v0/q2 [8]),
    .B1(\v0/z6/_018_ ),
    .Y(\v0/z6/_022_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z6/_165_  (.A(\v0/z6/_021_ ),
    .B(\v0/z6/_022_ ),
    .Y(\v0/q5 [9]));
 sky130_fd_sc_hd__nand2_1 \v0/z6/_166_  (.A(\v0/q3 [2]),
    .B(\v0/q2 [10]),
    .Y(\v0/z6/_023_ ));
 sky130_fd_sc_hd__xor2_1 \v0/z6/_167_  (.A(\v0/q3 [2]),
    .B(\v0/q2 [10]),
    .X(\v0/z6/_024_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z6/_168_  (.A(\v0/z6/_014_ ),
    .B(\v0/z6/_020_ ),
    .Y(\v0/z6/_025_ ));
 sky130_fd_sc_hd__o21ai_0 \v0/z6/_169_  (.A1(\v0/z6/_018_ ),
    .A2(\v0/z6/_025_ ),
    .B1(\v0/z6/_019_ ),
    .Y(\v0/z6/_026_ ));
 sky130_fd_sc_hd__o211ai_1 \v0/z6/_170_  (.A1(\v0/z6/_018_ ),
    .A2(\v0/z6/_025_ ),
    .B1(\v0/z6/_024_ ),
    .C1(\v0/z6/_019_ ),
    .Y(\v0/z6/_027_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z6/_171_  (.A(\v0/z6/_024_ ),
    .B(\v0/z6/_026_ ),
    .Y(\v0/q5 [10]));
 sky130_fd_sc_hd__nor2_1 \v0/z6/_172_  (.A(\v0/q3 [3]),
    .B(\v0/q2 [11]),
    .Y(\v0/z6/_028_ ));
 sky130_fd_sc_hd__lpflow_inputiso1p_1 \v0/z6/_173_  (.A(\v0/q3 [3]),
    .SLEEP(\v0/q2 [11]),
    .X(\v0/z6/_029_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z6/_174_  (.A(\v0/q3 [3]),
    .B(\v0/q2 [11]),
    .Y(\v0/z6/_030_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z6/_175_  (.A(\v0/z6/_029_ ),
    .B(\v0/z6/_030_ ),
    .Y(\v0/z6/_031_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z6/_176_  (.A(\v0/z6/_023_ ),
    .B(\v0/z6/_027_ ),
    .Y(\v0/z6/_032_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z6/_177_  (.A(\v0/z6/_031_ ),
    .B(\v0/z6/_032_ ),
    .Y(\v0/q5 [11]));
 sky130_fd_sc_hd__nand2_1 \v0/z6/_178_  (.A(\v0/q3 [4]),
    .B(\v0/q2 [12]),
    .Y(\v0/z6/_033_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z6/_179_  (.A(\v0/q3 [4]),
    .B(\v0/q2 [12]),
    .Y(\v0/z6/_034_ ));
 sky130_fd_sc_hd__and2_0 \v0/z6/_180_  (.A(\v0/z6/_023_ ),
    .B(\v0/z6/_030_ ),
    .X(\v0/z6/_035_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z6/_181_  (.A(\v0/z6/_027_ ),
    .B(\v0/z6/_035_ ),
    .Y(\v0/z6/_036_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z6/_182_  (.A(\v0/z6/_029_ ),
    .B(\v0/z6/_036_ ),
    .Y(\v0/z6/_037_ ));
 sky130_fd_sc_hd__a211oi_1 \v0/z6/_183_  (.A1(\v0/z6/_027_ ),
    .A2(\v0/z6/_035_ ),
    .B1(\v0/z6/_034_ ),
    .C1(\v0/z6/_028_ ),
    .Y(\v0/z6/_038_ ));
 sky130_fd_sc_hd__xor2_1 \v0/z6/_184_  (.A(\v0/z6/_034_ ),
    .B(\v0/z6/_037_ ),
    .X(\v0/q5 [12]));
 sky130_fd_sc_hd__lpflow_inputiso1p_1 \v0/z6/_185_  (.A(\v0/q3 [5]),
    .SLEEP(\v0/q2 [13]),
    .X(\v0/z6/_039_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z6/_186_  (.A(\v0/q3 [5]),
    .B(\v0/q2 [13]),
    .Y(\v0/z6/_040_ ));
 sky130_fd_sc_hd__and2_0 \v0/z6/_187_  (.A(\v0/z6/_039_ ),
    .B(\v0/z6/_040_ ),
    .X(\v0/z6/_041_ ));
 sky130_fd_sc_hd__a21oi_1 \v0/z6/_188_  (.A1(\v0/q3 [4]),
    .A2(\v0/q2 [12]),
    .B1(\v0/z6/_038_ ),
    .Y(\v0/z6/_042_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z6/_189_  (.A(\v0/z6/_041_ ),
    .B(\v0/z6/_042_ ),
    .Y(\v0/q5 [13]));
 sky130_fd_sc_hd__nand2_1 \v0/z6/_190_  (.A(\v0/q3 [6]),
    .B(\v0/q2 [14]),
    .Y(\v0/z6/_043_ ));
 sky130_fd_sc_hd__xor2_1 \v0/z6/_191_  (.A(\v0/q3 [6]),
    .B(\v0/q2 [14]),
    .X(\v0/z6/_044_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z6/_192_  (.A(\v0/z6/_033_ ),
    .B(\v0/z6/_040_ ),
    .Y(\v0/z6/_045_ ));
 sky130_fd_sc_hd__o21ai_0 \v0/z6/_193_  (.A1(\v0/z6/_038_ ),
    .A2(\v0/z6/_045_ ),
    .B1(\v0/z6/_039_ ),
    .Y(\v0/z6/_046_ ));
 sky130_fd_sc_hd__o211ai_1 \v0/z6/_194_  (.A1(\v0/z6/_038_ ),
    .A2(\v0/z6/_045_ ),
    .B1(\v0/z6/_044_ ),
    .C1(\v0/z6/_039_ ),
    .Y(\v0/z6/_047_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z6/_195_  (.A(\v0/z6/_044_ ),
    .B(\v0/z6/_046_ ),
    .Y(\v0/q5 [14]));
 sky130_fd_sc_hd__nand2_1 \v0/z6/_196_  (.A(\v0/q3 [7]),
    .B(\v0/q2 [15]),
    .Y(\v0/z6/_048_ ));
 sky130_fd_sc_hd__clkinv_1 \v0/z6/_197_  (.A(\v0/z6/_048_ ),
    .Y(\v0/z6/_049_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z6/_198_  (.A(\v0/q3 [7]),
    .B(\v0/q2 [15]),
    .Y(\v0/z6/_050_ ));
 sky130_fd_sc_hd__a21oi_1 \v0/z6/_199_  (.A1(\v0/z6/_043_ ),
    .A2(\v0/z6/_047_ ),
    .B1(\v0/z6/_050_ ),
    .Y(\v0/z6/_051_ ));
 sky130_fd_sc_hd__nand3_1 \v0/z6/_200_  (.A(\v0/z6/_043_ ),
    .B(\v0/z6/_047_ ),
    .C(\v0/z6/_050_ ),
    .Y(\v0/z6/_052_ ));
 sky130_fd_sc_hd__nor2b_1 \v0/z6/_201_  (.A(\v0/z6/_051_ ),
    .B_N(\v0/z6/_052_ ),
    .Y(\v0/q5 [15]));
 sky130_fd_sc_hd__lpflow_inputiso1p_1 \v0/z6/_202_  (.A(\v0/q3 [8]),
    .SLEEP(\v0/_09_ ),
    .X(\v0/z6/_053_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z6/_203_  (.A(\v0/q3 [8]),
    .B(\v0/_09_ ),
    .Y(\v0/z6/_054_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z6/_204_  (.A(\v0/z6/_053_ ),
    .B(\v0/z6/_054_ ),
    .Y(\v0/z6/_055_ ));
 sky130_fd_sc_hd__nor2_1 \v0/z6/_205_  (.A(\v0/z6/_049_ ),
    .B(\v0/z6/_051_ ),
    .Y(\v0/z6/_056_ ));
 sky130_fd_sc_hd__o21bai_1 \v0/z6/_206_  (.A1(\v0/z6/_049_ ),
    .A2(\v0/z6/_051_ ),
    .B1_N(\v0/z6/_055_ ),
    .Y(\v0/z6/_057_ ));
 sky130_fd_sc_hd__xor2_1 \v0/z6/_207_  (.A(\v0/z6/_055_ ),
    .B(\v0/z6/_056_ ),
    .X(\v0/q5 [16]));
 sky130_fd_sc_hd__nor2_1 \v0/z6/_208_  (.A(\v0/q3 [9]),
    .B(\v0/_10_ ),
    .Y(\v0/z6/_058_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z6/_209_  (.A(\v0/q3 [9]),
    .B(\v0/_10_ ),
    .Y(\v0/z6/_059_ ));
 sky130_fd_sc_hd__nor2b_1 \v0/z6/_210_  (.A(\v0/z6/_058_ ),
    .B_N(\v0/z6/_059_ ),
    .Y(\v0/z6/_060_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z6/_211_  (.A(\v0/z6/_048_ ),
    .B(\v0/z6/_054_ ),
    .Y(\v0/z6/_061_ ));
 sky130_fd_sc_hd__o21ai_0 \v0/z6/_212_  (.A1(\v0/z6/_051_ ),
    .A2(\v0/z6/_061_ ),
    .B1(\v0/z6/_053_ ),
    .Y(\v0/z6/_062_ ));
 sky130_fd_sc_hd__o211ai_1 \v0/z6/_213_  (.A1(\v0/z6/_051_ ),
    .A2(\v0/z6/_061_ ),
    .B1(\v0/z6/_060_ ),
    .C1(\v0/z6/_053_ ),
    .Y(\v0/z6/_063_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z6/_214_  (.A(\v0/z6/_060_ ),
    .B(\v0/z6/_062_ ),
    .Y(\v0/q5 [17]));
 sky130_fd_sc_hd__nor2_1 \v0/z6/_215_  (.A(\v0/q3 [10]),
    .B(\v0/_11_ ),
    .Y(\v0/z6/_064_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z6/_216_  (.A(\v0/q3 [10]),
    .B(\v0/_11_ ),
    .Y(\v0/z6/_065_ ));
 sky130_fd_sc_hd__nand2b_1 \v0/z6/_217_  (.A_N(\v0/z6/_064_ ),
    .B(\v0/z6/_065_ ),
    .Y(\v0/z6/_066_ ));
 sky130_fd_sc_hd__a31oi_1 \v0/z6/_218_  (.A1(\v0/z6/_054_ ),
    .A2(\v0/z6/_057_ ),
    .A3(\v0/z6/_059_ ),
    .B1(\v0/z6/_058_ ),
    .Y(\v0/z6/_067_ ));
 sky130_fd_sc_hd__a311o_1 \v0/z6/_219_  (.A1(\v0/z6/_054_ ),
    .A2(\v0/z6/_057_ ),
    .A3(\v0/z6/_059_ ),
    .B1(\v0/z6/_066_ ),
    .C1(\v0/z6/_058_ ),
    .X(\v0/z6/_068_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z6/_220_  (.A(\v0/z6/_066_ ),
    .B(\v0/z6/_067_ ),
    .Y(\v0/q5 [18]));
 sky130_fd_sc_hd__nor2_1 \v0/z6/_221_  (.A(\v0/q3 [11]),
    .B(\v0/_12_ ),
    .Y(\v0/z6/_069_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z6/_222_  (.A(\v0/q3 [11]),
    .B(\v0/_12_ ),
    .Y(\v0/z6/_070_ ));
 sky130_fd_sc_hd__nand2b_1 \v0/z6/_223_  (.A_N(\v0/z6/_069_ ),
    .B(\v0/z6/_070_ ),
    .Y(\v0/z6/_071_ ));
 sky130_fd_sc_hd__a31oi_1 \v0/z6/_224_  (.A1(\v0/z6/_059_ ),
    .A2(\v0/z6/_063_ ),
    .A3(\v0/z6/_065_ ),
    .B1(\v0/z6/_064_ ),
    .Y(\v0/z6/_072_ ));
 sky130_fd_sc_hd__a311oi_1 \v0/z6/_225_  (.A1(\v0/z6/_059_ ),
    .A2(\v0/z6/_063_ ),
    .A3(\v0/z6/_065_ ),
    .B1(\v0/z6/_071_ ),
    .C1(\v0/z6/_064_ ),
    .Y(\v0/z6/_073_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z6/_226_  (.A(\v0/z6/_071_ ),
    .B(\v0/z6/_072_ ),
    .Y(\v0/q5 [19]));
 sky130_fd_sc_hd__nand2_1 \v0/z6/_227_  (.A(\v0/q3 [12]),
    .B(\v0/_13_ ),
    .Y(\v0/z6/_074_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z6/_228_  (.A(\v0/q3 [12]),
    .B(\v0/_13_ ),
    .Y(\v0/z6/_075_ ));
 sky130_fd_sc_hd__a31oi_1 \v0/z6/_229_  (.A1(\v0/z6/_065_ ),
    .A2(\v0/z6/_068_ ),
    .A3(\v0/z6/_070_ ),
    .B1(\v0/z6/_069_ ),
    .Y(\v0/z6/_076_ ));
 sky130_fd_sc_hd__a311o_1 \v0/z6/_230_  (.A1(\v0/z6/_065_ ),
    .A2(\v0/z6/_068_ ),
    .A3(\v0/z6/_070_ ),
    .B1(\v0/z6/_075_ ),
    .C1(\v0/z6/_069_ ),
    .X(\v0/z6/_077_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z6/_231_  (.A(\v0/z6/_075_ ),
    .B(\v0/z6/_076_ ),
    .Y(\v0/q5 [20]));
 sky130_fd_sc_hd__nor2_1 \v0/z6/_232_  (.A(\v0/q3 [13]),
    .B(\v0/_14_ ),
    .Y(\v0/z6/_078_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z6/_233_  (.A(\v0/q3 [13]),
    .B(\v0/_14_ ),
    .Y(\v0/z6/_079_ ));
 sky130_fd_sc_hd__nor2b_1 \v0/z6/_234_  (.A(\v0/z6/_078_ ),
    .B_N(\v0/z6/_079_ ),
    .Y(\v0/z6/_080_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z6/_235_  (.A(\v0/z6/_070_ ),
    .B(\v0/z6/_074_ ),
    .Y(\v0/z6/_081_ ));
 sky130_fd_sc_hd__o22ai_1 \v0/z6/_236_  (.A1(\v0/q3 [12]),
    .A2(\v0/_13_ ),
    .B1(\v0/z6/_073_ ),
    .B2(\v0/z6/_081_ ),
    .Y(\v0/z6/_082_ ));
 sky130_fd_sc_hd__o221ai_1 \v0/z6/_237_  (.A1(\v0/q3 [12]),
    .A2(\v0/_13_ ),
    .B1(\v0/z6/_073_ ),
    .B2(\v0/z6/_081_ ),
    .C1(\v0/z6/_080_ ),
    .Y(\v0/z6/_083_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z6/_238_  (.A(\v0/z6/_080_ ),
    .B(\v0/z6/_082_ ),
    .Y(\v0/q5 [21]));
 sky130_fd_sc_hd__nor2_1 \v0/z6/_239_  (.A(\v0/q3 [14]),
    .B(\v0/_15_ ),
    .Y(\v0/z6/_084_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z6/_240_  (.A(\v0/q3 [14]),
    .B(\v0/_15_ ),
    .Y(\v0/z6/_085_ ));
 sky130_fd_sc_hd__nand2b_1 \v0/z6/_241_  (.A_N(\v0/z6/_084_ ),
    .B(\v0/z6/_085_ ),
    .Y(\v0/z6/_086_ ));
 sky130_fd_sc_hd__a31oi_1 \v0/z6/_242_  (.A1(\v0/z6/_074_ ),
    .A2(\v0/z6/_077_ ),
    .A3(\v0/z6/_079_ ),
    .B1(\v0/z6/_078_ ),
    .Y(\v0/z6/_087_ ));
 sky130_fd_sc_hd__a311o_1 \v0/z6/_243_  (.A1(\v0/z6/_074_ ),
    .A2(\v0/z6/_077_ ),
    .A3(\v0/z6/_079_ ),
    .B1(\v0/z6/_086_ ),
    .C1(\v0/z6/_078_ ),
    .X(\v0/z6/_088_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z6/_244_  (.A(\v0/z6/_086_ ),
    .B(\v0/z6/_087_ ),
    .Y(\v0/q5 [22]));
 sky130_fd_sc_hd__nor2_1 \v0/z6/_245_  (.A(\v0/q3 [15]),
    .B(\v0/_16_ ),
    .Y(\v0/z6/_089_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z6/_246_  (.A(\v0/q3 [15]),
    .B(\v0/_16_ ),
    .Y(\v0/z6/_090_ ));
 sky130_fd_sc_hd__nand2b_1 \v0/z6/_247_  (.A_N(\v0/z6/_089_ ),
    .B(\v0/z6/_090_ ),
    .Y(\v0/z6/_091_ ));
 sky130_fd_sc_hd__a31oi_1 \v0/z6/_248_  (.A1(\v0/z6/_079_ ),
    .A2(\v0/z6/_083_ ),
    .A3(\v0/z6/_085_ ),
    .B1(\v0/z6/_084_ ),
    .Y(\v0/z6/_092_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z6/_249_  (.A(\v0/z6/_091_ ),
    .B(\v0/z6/_092_ ),
    .Y(\v0/q5 [23]));
 sky130_fd_sc_hd__a31oi_1 \v0/z6/_250_  (.A1(\v0/z6/_085_ ),
    .A2(\v0/z6/_088_ ),
    .A3(\v0/z6/_090_ ),
    .B1(\v0/z6/_089_ ),
    .Y(\v0/z6/Cout ));
 sky130_fd_sc_hd__xnor2_1 \v0/z7/_113_  (.A(\v0/q5 [0]),
    .B(\v0/q4 [0]),
    .Y(\v0/z7/_093_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z7/_114_  (.A(\v0/_34_ ),
    .B(\v0/z7/_093_ ),
    .Y(unsign[8]));
 sky130_fd_sc_hd__maj3_1 \v0/z7/_115_  (.A(\v0/q5 [0]),
    .B(\v0/q4 [0]),
    .C(\v0/_34_ ),
    .X(\v0/z7/_094_ ));
 sky130_fd_sc_hd__lpflow_inputiso1p_1 \v0/z7/_116_  (.A(\v0/q5 [1]),
    .SLEEP(\v0/q4 [1]),
    .X(\v0/z7/_095_ ));
 sky130_fd_sc_hd__and2_0 \v0/z7/_117_  (.A(\v0/q5 [1]),
    .B(\v0/q4 [1]),
    .X(\v0/z7/_096_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z7/_118_  (.A(\v0/q5 [1]),
    .B(\v0/q4 [1]),
    .Y(\v0/z7/_097_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z7/_119_  (.A(\v0/z7/_095_ ),
    .B(\v0/z7/_097_ ),
    .Y(\v0/z7/_098_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z7/_120_  (.A(\v0/z7/_094_ ),
    .B(\v0/z7/_098_ ),
    .Y(unsign[9]));
 sky130_fd_sc_hd__nor2_1 \v0/z7/_121_  (.A(\v0/q5 [2]),
    .B(\v0/q4 [2]),
    .Y(\v0/z7/_099_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z7/_122_  (.A(\v0/q5 [2]),
    .B(\v0/q4 [2]),
    .Y(\v0/z7/_100_ ));
 sky130_fd_sc_hd__xor2_1 \v0/z7/_123_  (.A(\v0/q5 [2]),
    .B(\v0/q4 [2]),
    .X(\v0/z7/_101_ ));
 sky130_fd_sc_hd__o21ai_0 \v0/z7/_124_  (.A1(\v0/z7/_094_ ),
    .A2(\v0/z7/_096_ ),
    .B1(\v0/z7/_095_ ),
    .Y(\v0/z7/_102_ ));
 sky130_fd_sc_hd__o211a_1 \v0/z7/_125_  (.A1(\v0/z7/_094_ ),
    .A2(\v0/z7/_096_ ),
    .B1(\v0/z7/_101_ ),
    .C1(\v0/z7/_095_ ),
    .X(\v0/z7/_103_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z7/_126_  (.A(\v0/z7/_101_ ),
    .B(\v0/z7/_102_ ),
    .Y(unsign[10]));
 sky130_fd_sc_hd__nand2_1 \v0/z7/_127_  (.A(\v0/q5 [3]),
    .B(\v0/q4 [3]),
    .Y(\v0/z7/_104_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z7/_128_  (.A(\v0/q5 [3]),
    .B(\v0/q4 [3]),
    .Y(\v0/z7/_105_ ));
 sky130_fd_sc_hd__o21ai_0 \v0/z7/_129_  (.A1(\v0/z7/_099_ ),
    .A2(\v0/z7/_102_ ),
    .B1(\v0/z7/_100_ ),
    .Y(\v0/z7/_106_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z7/_130_  (.A(\v0/z7/_105_ ),
    .B(\v0/z7/_106_ ),
    .Y(unsign[11]));
 sky130_fd_sc_hd__lpflow_inputiso1p_1 \v0/z7/_131_  (.A(\v0/q5 [4]),
    .SLEEP(\v0/q4 [4]),
    .X(\v0/z7/_107_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z7/_132_  (.A(\v0/q5 [4]),
    .B(\v0/q4 [4]),
    .Y(\v0/z7/_108_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z7/_133_  (.A(\v0/z7/_107_ ),
    .B(\v0/z7/_108_ ),
    .Y(\v0/z7/_109_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z7/_134_  (.A(\v0/z7/_100_ ),
    .B(\v0/z7/_104_ ),
    .Y(\v0/z7/_110_ ));
 sky130_fd_sc_hd__o22a_1 \v0/z7/_135_  (.A1(\v0/q5 [3]),
    .A2(\v0/q4 [3]),
    .B1(\v0/z7/_103_ ),
    .B2(\v0/z7/_110_ ),
    .X(\v0/z7/_111_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z7/_136_  (.A(\v0/z7/_109_ ),
    .B(\v0/z7/_111_ ),
    .Y(unsign[12]));
 sky130_fd_sc_hd__nor2_1 \v0/z7/_137_  (.A(\v0/q5 [5]),
    .B(\v0/q4 [5]),
    .Y(\v0/z7/_112_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z7/_138_  (.A(\v0/q5 [5]),
    .B(\v0/q4 [5]),
    .Y(\v0/z7/_000_ ));
 sky130_fd_sc_hd__nand2b_1 \v0/z7/_139_  (.A_N(\v0/z7/_112_ ),
    .B(\v0/z7/_000_ ),
    .Y(\v0/z7/_001_ ));
 sky130_fd_sc_hd__o221ai_1 \v0/z7/_140_  (.A1(\v0/q5 [3]),
    .A2(\v0/q4 [3]),
    .B1(\v0/z7/_103_ ),
    .B2(\v0/z7/_110_ ),
    .C1(\v0/z7/_107_ ),
    .Y(\v0/z7/_002_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z7/_141_  (.A(\v0/z7/_108_ ),
    .B(\v0/z7/_002_ ),
    .Y(\v0/z7/_003_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z7/_142_  (.A(\v0/z7/_001_ ),
    .B(\v0/z7/_003_ ),
    .Y(unsign[13]));
 sky130_fd_sc_hd__nor2_1 \v0/z7/_143_  (.A(\v0/q5 [6]),
    .B(\v0/q4 [6]),
    .Y(\v0/z7/_004_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z7/_144_  (.A(\v0/q5 [6]),
    .B(\v0/q4 [6]),
    .Y(\v0/z7/_005_ ));
 sky130_fd_sc_hd__nor2b_1 \v0/z7/_145_  (.A(\v0/z7/_004_ ),
    .B_N(\v0/z7/_005_ ),
    .Y(\v0/z7/_006_ ));
 sky130_fd_sc_hd__clkinv_1 \v0/z7/_146_  (.A(\v0/z7/_006_ ),
    .Y(\v0/z7/_007_ ));
 sky130_fd_sc_hd__o21ai_0 \v0/z7/_147_  (.A1(\v0/q5 [5]),
    .A2(\v0/q4 [5]),
    .B1(\v0/z7/_003_ ),
    .Y(\v0/z7/_008_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z7/_148_  (.A(\v0/z7/_000_ ),
    .B(\v0/z7/_008_ ),
    .Y(\v0/z7/_009_ ));
 sky130_fd_sc_hd__a311o_1 \v0/z7/_149_  (.A1(\v0/z7/_108_ ),
    .A2(\v0/z7/_000_ ),
    .A3(\v0/z7/_002_ ),
    .B1(\v0/z7/_007_ ),
    .C1(\v0/z7/_112_ ),
    .X(\v0/z7/_010_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z7/_150_  (.A(\v0/z7/_007_ ),
    .B(\v0/z7/_009_ ),
    .Y(unsign[14]));
 sky130_fd_sc_hd__nor2_1 \v0/z7/_151_  (.A(\v0/q5 [7]),
    .B(\v0/q4 [7]),
    .Y(\v0/z7/_011_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z7/_152_  (.A(\v0/q5 [7]),
    .B(\v0/q4 [7]),
    .Y(\v0/z7/_012_ ));
 sky130_fd_sc_hd__a31oi_1 \v0/z7/_153_  (.A1(\v0/z7/_000_ ),
    .A2(\v0/z7/_005_ ),
    .A3(\v0/z7/_008_ ),
    .B1(\v0/z7/_004_ ),
    .Y(\v0/z7/_013_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z7/_154_  (.A(\v0/z7/_012_ ),
    .B(\v0/z7/_013_ ),
    .Y(unsign[15]));
 sky130_fd_sc_hd__nand2_1 \v0/z7/_155_  (.A(\v0/q5 [8]),
    .B(\v0/q4 [8]),
    .Y(\v0/z7/_014_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z7/_156_  (.A(\v0/q5 [8]),
    .B(\v0/q4 [8]),
    .Y(\v0/z7/_015_ ));
 sky130_fd_sc_hd__a22oi_1 \v0/z7/_157_  (.A1(\v0/q5 [6]),
    .A2(\v0/q4 [6]),
    .B1(\v0/q5 [7]),
    .B2(\v0/q4 [7]),
    .Y(\v0/z7/_016_ ));
 sky130_fd_sc_hd__a21oi_1 \v0/z7/_158_  (.A1(\v0/z7/_010_ ),
    .A2(\v0/z7/_016_ ),
    .B1(\v0/z7/_011_ ),
    .Y(\v0/z7/_017_ ));
 sky130_fd_sc_hd__a211oi_1 \v0/z7/_159_  (.A1(\v0/z7/_010_ ),
    .A2(\v0/z7/_016_ ),
    .B1(\v0/z7/_015_ ),
    .C1(\v0/z7/_011_ ),
    .Y(\v0/z7/_018_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z7/_160_  (.A(\v0/z7/_015_ ),
    .B(\v0/z7/_017_ ),
    .Y(unsign[16]));
 sky130_fd_sc_hd__lpflow_inputiso1p_1 \v0/z7/_161_  (.A(\v0/q5 [9]),
    .SLEEP(\v0/q4 [9]),
    .X(\v0/z7/_019_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z7/_162_  (.A(\v0/q5 [9]),
    .B(\v0/q4 [9]),
    .Y(\v0/z7/_020_ ));
 sky130_fd_sc_hd__and2_0 \v0/z7/_163_  (.A(\v0/z7/_019_ ),
    .B(\v0/z7/_020_ ),
    .X(\v0/z7/_021_ ));
 sky130_fd_sc_hd__a21oi_1 \v0/z7/_164_  (.A1(\v0/q5 [8]),
    .A2(\v0/q4 [8]),
    .B1(\v0/z7/_018_ ),
    .Y(\v0/z7/_022_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z7/_165_  (.A(\v0/z7/_021_ ),
    .B(\v0/z7/_022_ ),
    .Y(unsign[17]));
 sky130_fd_sc_hd__nand2_1 \v0/z7/_166_  (.A(\v0/q5 [10]),
    .B(\v0/q4 [10]),
    .Y(\v0/z7/_023_ ));
 sky130_fd_sc_hd__xor2_1 \v0/z7/_167_  (.A(\v0/q5 [10]),
    .B(\v0/q4 [10]),
    .X(\v0/z7/_024_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z7/_168_  (.A(\v0/z7/_014_ ),
    .B(\v0/z7/_020_ ),
    .Y(\v0/z7/_025_ ));
 sky130_fd_sc_hd__o21ai_0 \v0/z7/_169_  (.A1(\v0/z7/_018_ ),
    .A2(\v0/z7/_025_ ),
    .B1(\v0/z7/_019_ ),
    .Y(\v0/z7/_026_ ));
 sky130_fd_sc_hd__o211ai_1 \v0/z7/_170_  (.A1(\v0/z7/_018_ ),
    .A2(\v0/z7/_025_ ),
    .B1(\v0/z7/_024_ ),
    .C1(\v0/z7/_019_ ),
    .Y(\v0/z7/_027_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z7/_171_  (.A(\v0/z7/_024_ ),
    .B(\v0/z7/_026_ ),
    .Y(unsign[18]));
 sky130_fd_sc_hd__nor2_1 \v0/z7/_172_  (.A(\v0/q5 [11]),
    .B(\v0/q4 [11]),
    .Y(\v0/z7/_028_ ));
 sky130_fd_sc_hd__lpflow_inputiso1p_1 \v0/z7/_173_  (.A(\v0/q5 [11]),
    .SLEEP(\v0/q4 [11]),
    .X(\v0/z7/_029_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z7/_174_  (.A(\v0/q5 [11]),
    .B(\v0/q4 [11]),
    .Y(\v0/z7/_030_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z7/_175_  (.A(\v0/z7/_029_ ),
    .B(\v0/z7/_030_ ),
    .Y(\v0/z7/_031_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z7/_176_  (.A(\v0/z7/_023_ ),
    .B(\v0/z7/_027_ ),
    .Y(\v0/z7/_032_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z7/_177_  (.A(\v0/z7/_031_ ),
    .B(\v0/z7/_032_ ),
    .Y(unsign[19]));
 sky130_fd_sc_hd__nand2_1 \v0/z7/_178_  (.A(\v0/q5 [12]),
    .B(\v0/q4 [12]),
    .Y(\v0/z7/_033_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z7/_179_  (.A(\v0/q5 [12]),
    .B(\v0/q4 [12]),
    .Y(\v0/z7/_034_ ));
 sky130_fd_sc_hd__and2_0 \v0/z7/_180_  (.A(\v0/z7/_023_ ),
    .B(\v0/z7/_030_ ),
    .X(\v0/z7/_035_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z7/_181_  (.A(\v0/z7/_027_ ),
    .B(\v0/z7/_035_ ),
    .Y(\v0/z7/_036_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z7/_182_  (.A(\v0/z7/_029_ ),
    .B(\v0/z7/_036_ ),
    .Y(\v0/z7/_037_ ));
 sky130_fd_sc_hd__a211oi_1 \v0/z7/_183_  (.A1(\v0/z7/_027_ ),
    .A2(\v0/z7/_035_ ),
    .B1(\v0/z7/_034_ ),
    .C1(\v0/z7/_028_ ),
    .Y(\v0/z7/_038_ ));
 sky130_fd_sc_hd__xor2_1 \v0/z7/_184_  (.A(\v0/z7/_034_ ),
    .B(\v0/z7/_037_ ),
    .X(unsign[20]));
 sky130_fd_sc_hd__lpflow_inputiso1p_1 \v0/z7/_185_  (.A(\v0/q5 [13]),
    .SLEEP(\v0/q4 [13]),
    .X(\v0/z7/_039_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z7/_186_  (.A(\v0/q5 [13]),
    .B(\v0/q4 [13]),
    .Y(\v0/z7/_040_ ));
 sky130_fd_sc_hd__and2_0 \v0/z7/_187_  (.A(\v0/z7/_039_ ),
    .B(\v0/z7/_040_ ),
    .X(\v0/z7/_041_ ));
 sky130_fd_sc_hd__a21oi_1 \v0/z7/_188_  (.A1(\v0/q5 [12]),
    .A2(\v0/q4 [12]),
    .B1(\v0/z7/_038_ ),
    .Y(\v0/z7/_042_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z7/_189_  (.A(\v0/z7/_041_ ),
    .B(\v0/z7/_042_ ),
    .Y(unsign[21]));
 sky130_fd_sc_hd__nand2_1 \v0/z7/_190_  (.A(\v0/q5 [14]),
    .B(\v0/q4 [14]),
    .Y(\v0/z7/_043_ ));
 sky130_fd_sc_hd__xor2_1 \v0/z7/_191_  (.A(\v0/q5 [14]),
    .B(\v0/q4 [14]),
    .X(\v0/z7/_044_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z7/_192_  (.A(\v0/z7/_033_ ),
    .B(\v0/z7/_040_ ),
    .Y(\v0/z7/_045_ ));
 sky130_fd_sc_hd__o21ai_0 \v0/z7/_193_  (.A1(\v0/z7/_038_ ),
    .A2(\v0/z7/_045_ ),
    .B1(\v0/z7/_039_ ),
    .Y(\v0/z7/_046_ ));
 sky130_fd_sc_hd__o211ai_1 \v0/z7/_194_  (.A1(\v0/z7/_038_ ),
    .A2(\v0/z7/_045_ ),
    .B1(\v0/z7/_044_ ),
    .C1(\v0/z7/_039_ ),
    .Y(\v0/z7/_047_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z7/_195_  (.A(\v0/z7/_044_ ),
    .B(\v0/z7/_046_ ),
    .Y(unsign[22]));
 sky130_fd_sc_hd__nand2_1 \v0/z7/_196_  (.A(\v0/q5 [15]),
    .B(\v0/q4 [15]),
    .Y(\v0/z7/_048_ ));
 sky130_fd_sc_hd__clkinv_1 \v0/z7/_197_  (.A(\v0/z7/_048_ ),
    .Y(\v0/z7/_049_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z7/_198_  (.A(\v0/q5 [15]),
    .B(\v0/q4 [15]),
    .Y(\v0/z7/_050_ ));
 sky130_fd_sc_hd__a21oi_1 \v0/z7/_199_  (.A1(\v0/z7/_043_ ),
    .A2(\v0/z7/_047_ ),
    .B1(\v0/z7/_050_ ),
    .Y(\v0/z7/_051_ ));
 sky130_fd_sc_hd__nand3_1 \v0/z7/_200_  (.A(\v0/z7/_043_ ),
    .B(\v0/z7/_047_ ),
    .C(\v0/z7/_050_ ),
    .Y(\v0/z7/_052_ ));
 sky130_fd_sc_hd__nor2b_1 \v0/z7/_201_  (.A(\v0/z7/_051_ ),
    .B_N(\v0/z7/_052_ ),
    .Y(unsign[23]));
 sky130_fd_sc_hd__lpflow_inputiso1p_1 \v0/z7/_202_  (.A(\v0/q5 [16]),
    .SLEEP(\v0/_26_ ),
    .X(\v0/z7/_053_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z7/_203_  (.A(\v0/q5 [16]),
    .B(\v0/_26_ ),
    .Y(\v0/z7/_054_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z7/_204_  (.A(\v0/z7/_053_ ),
    .B(\v0/z7/_054_ ),
    .Y(\v0/z7/_055_ ));
 sky130_fd_sc_hd__nor2_1 \v0/z7/_205_  (.A(\v0/z7/_049_ ),
    .B(\v0/z7/_051_ ),
    .Y(\v0/z7/_056_ ));
 sky130_fd_sc_hd__o21bai_1 \v0/z7/_206_  (.A1(\v0/z7/_049_ ),
    .A2(\v0/z7/_051_ ),
    .B1_N(\v0/z7/_055_ ),
    .Y(\v0/z7/_057_ ));
 sky130_fd_sc_hd__xor2_1 \v0/z7/_207_  (.A(\v0/z7/_055_ ),
    .B(\v0/z7/_056_ ),
    .X(unsign[24]));
 sky130_fd_sc_hd__nor2_1 \v0/z7/_208_  (.A(\v0/q5 [17]),
    .B(\v0/_27_ ),
    .Y(\v0/z7/_058_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z7/_209_  (.A(\v0/q5 [17]),
    .B(\v0/_27_ ),
    .Y(\v0/z7/_059_ ));
 sky130_fd_sc_hd__nor2b_1 \v0/z7/_210_  (.A(\v0/z7/_058_ ),
    .B_N(\v0/z7/_059_ ),
    .Y(\v0/z7/_060_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z7/_211_  (.A(\v0/z7/_048_ ),
    .B(\v0/z7/_054_ ),
    .Y(\v0/z7/_061_ ));
 sky130_fd_sc_hd__o21ai_0 \v0/z7/_212_  (.A1(\v0/z7/_051_ ),
    .A2(\v0/z7/_061_ ),
    .B1(\v0/z7/_053_ ),
    .Y(\v0/z7/_062_ ));
 sky130_fd_sc_hd__o211ai_1 \v0/z7/_213_  (.A1(\v0/z7/_051_ ),
    .A2(\v0/z7/_061_ ),
    .B1(\v0/z7/_060_ ),
    .C1(\v0/z7/_053_ ),
    .Y(\v0/z7/_063_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z7/_214_  (.A(\v0/z7/_060_ ),
    .B(\v0/z7/_062_ ),
    .Y(unsign[25]));
 sky130_fd_sc_hd__nor2_1 \v0/z7/_215_  (.A(\v0/q5 [18]),
    .B(\v0/_28_ ),
    .Y(\v0/z7/_064_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z7/_216_  (.A(\v0/q5 [18]),
    .B(\v0/_28_ ),
    .Y(\v0/z7/_065_ ));
 sky130_fd_sc_hd__nand2b_1 \v0/z7/_217_  (.A_N(\v0/z7/_064_ ),
    .B(\v0/z7/_065_ ),
    .Y(\v0/z7/_066_ ));
 sky130_fd_sc_hd__a31oi_1 \v0/z7/_218_  (.A1(\v0/z7/_054_ ),
    .A2(\v0/z7/_057_ ),
    .A3(\v0/z7/_059_ ),
    .B1(\v0/z7/_058_ ),
    .Y(\v0/z7/_067_ ));
 sky130_fd_sc_hd__a311o_1 \v0/z7/_219_  (.A1(\v0/z7/_054_ ),
    .A2(\v0/z7/_057_ ),
    .A3(\v0/z7/_059_ ),
    .B1(\v0/z7/_066_ ),
    .C1(\v0/z7/_058_ ),
    .X(\v0/z7/_068_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z7/_220_  (.A(\v0/z7/_066_ ),
    .B(\v0/z7/_067_ ),
    .Y(unsign[26]));
 sky130_fd_sc_hd__nor2_1 \v0/z7/_221_  (.A(\v0/q5 [19]),
    .B(\v0/_29_ ),
    .Y(\v0/z7/_069_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z7/_222_  (.A(\v0/q5 [19]),
    .B(\v0/_29_ ),
    .Y(\v0/z7/_070_ ));
 sky130_fd_sc_hd__nand2b_1 \v0/z7/_223_  (.A_N(\v0/z7/_069_ ),
    .B(\v0/z7/_070_ ),
    .Y(\v0/z7/_071_ ));
 sky130_fd_sc_hd__a31oi_1 \v0/z7/_224_  (.A1(\v0/z7/_059_ ),
    .A2(\v0/z7/_063_ ),
    .A3(\v0/z7/_065_ ),
    .B1(\v0/z7/_064_ ),
    .Y(\v0/z7/_072_ ));
 sky130_fd_sc_hd__a311oi_1 \v0/z7/_225_  (.A1(\v0/z7/_059_ ),
    .A2(\v0/z7/_063_ ),
    .A3(\v0/z7/_065_ ),
    .B1(\v0/z7/_071_ ),
    .C1(\v0/z7/_064_ ),
    .Y(\v0/z7/_073_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z7/_226_  (.A(\v0/z7/_071_ ),
    .B(\v0/z7/_072_ ),
    .Y(unsign[27]));
 sky130_fd_sc_hd__nand2_1 \v0/z7/_227_  (.A(\v0/q5 [20]),
    .B(\v0/_30_ ),
    .Y(\v0/z7/_074_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z7/_228_  (.A(\v0/q5 [20]),
    .B(\v0/_30_ ),
    .Y(\v0/z7/_075_ ));
 sky130_fd_sc_hd__a31oi_1 \v0/z7/_229_  (.A1(\v0/z7/_065_ ),
    .A2(\v0/z7/_068_ ),
    .A3(\v0/z7/_070_ ),
    .B1(\v0/z7/_069_ ),
    .Y(\v0/z7/_076_ ));
 sky130_fd_sc_hd__a311o_1 \v0/z7/_230_  (.A1(\v0/z7/_065_ ),
    .A2(\v0/z7/_068_ ),
    .A3(\v0/z7/_070_ ),
    .B1(\v0/z7/_075_ ),
    .C1(\v0/z7/_069_ ),
    .X(\v0/z7/_077_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z7/_231_  (.A(\v0/z7/_075_ ),
    .B(\v0/z7/_076_ ),
    .Y(unsign[28]));
 sky130_fd_sc_hd__nor2_1 \v0/z7/_232_  (.A(\v0/q5 [21]),
    .B(\v0/_31_ ),
    .Y(\v0/z7/_078_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z7/_233_  (.A(\v0/q5 [21]),
    .B(\v0/_31_ ),
    .Y(\v0/z7/_079_ ));
 sky130_fd_sc_hd__nor2b_1 \v0/z7/_234_  (.A(\v0/z7/_078_ ),
    .B_N(\v0/z7/_079_ ),
    .Y(\v0/z7/_080_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z7/_235_  (.A(\v0/z7/_070_ ),
    .B(\v0/z7/_074_ ),
    .Y(\v0/z7/_081_ ));
 sky130_fd_sc_hd__o22ai_1 \v0/z7/_236_  (.A1(\v0/q5 [20]),
    .A2(\v0/_30_ ),
    .B1(\v0/z7/_073_ ),
    .B2(\v0/z7/_081_ ),
    .Y(\v0/z7/_082_ ));
 sky130_fd_sc_hd__o221ai_1 \v0/z7/_237_  (.A1(\v0/q5 [20]),
    .A2(\v0/_30_ ),
    .B1(\v0/z7/_073_ ),
    .B2(\v0/z7/_081_ ),
    .C1(\v0/z7/_080_ ),
    .Y(\v0/z7/_083_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z7/_238_  (.A(\v0/z7/_080_ ),
    .B(\v0/z7/_082_ ),
    .Y(unsign[29]));
 sky130_fd_sc_hd__nor2_1 \v0/z7/_239_  (.A(\v0/q5 [22]),
    .B(\v0/_32_ ),
    .Y(\v0/z7/_084_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z7/_240_  (.A(\v0/q5 [22]),
    .B(\v0/_32_ ),
    .Y(\v0/z7/_085_ ));
 sky130_fd_sc_hd__nand2b_1 \v0/z7/_241_  (.A_N(\v0/z7/_084_ ),
    .B(\v0/z7/_085_ ),
    .Y(\v0/z7/_086_ ));
 sky130_fd_sc_hd__a31oi_1 \v0/z7/_242_  (.A1(\v0/z7/_074_ ),
    .A2(\v0/z7/_077_ ),
    .A3(\v0/z7/_079_ ),
    .B1(\v0/z7/_078_ ),
    .Y(\v0/z7/_087_ ));
 sky130_fd_sc_hd__a311o_1 \v0/z7/_243_  (.A1(\v0/z7/_074_ ),
    .A2(\v0/z7/_077_ ),
    .A3(\v0/z7/_079_ ),
    .B1(\v0/z7/_086_ ),
    .C1(\v0/z7/_078_ ),
    .X(\v0/z7/_088_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z7/_244_  (.A(\v0/z7/_086_ ),
    .B(\v0/z7/_087_ ),
    .Y(unsign[30]));
 sky130_fd_sc_hd__nor2_1 \v0/z7/_245_  (.A(\v0/q5 [23]),
    .B(\v0/_33_ ),
    .Y(\v0/z7/_089_ ));
 sky130_fd_sc_hd__nand2_1 \v0/z7/_246_  (.A(\v0/q5 [23]),
    .B(\v0/_33_ ),
    .Y(\v0/z7/_090_ ));
 sky130_fd_sc_hd__nand2b_1 \v0/z7/_247_  (.A_N(\v0/z7/_089_ ),
    .B(\v0/z7/_090_ ),
    .Y(\v0/z7/_091_ ));
 sky130_fd_sc_hd__a31oi_1 \v0/z7/_248_  (.A1(\v0/z7/_079_ ),
    .A2(\v0/z7/_083_ ),
    .A3(\v0/z7/_085_ ),
    .B1(\v0/z7/_084_ ),
    .Y(\v0/z7/_092_ ));
 sky130_fd_sc_hd__xnor2_1 \v0/z7/_249_  (.A(\v0/z7/_091_ ),
    .B(\v0/z7/_092_ ),
    .Y(unsign[31]));
 sky130_fd_sc_hd__a31oi_1 \v0/z7/_250_  (.A1(\v0/z7/_085_ ),
    .A2(\v0/z7/_088_ ),
    .A3(\v0/z7/_090_ ),
    .B1(\v0/z7/_089_ ),
    .Y(\v0/z7/Cout ));
endmodule
